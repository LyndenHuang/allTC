VERSION 5.8 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 4000 ;
END UNITS

MANUFACTURINGGRID 0.0005 ;

PROPERTYDEFINITIONS
  MACRO write_qor_data STRING ;
  MACRO port_placement_export_file STRING ;
  MACRO sqs_step STRING ;
  MACRO rm_lib_type STRING ;
END PROPERTYDEFINITIONS

LAYER bsb
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 80 ;
  WIDTH 32 ;
  PROPERTY LEF58_WIDTH "WIDTH 32 WRONGDIRECTION ;" ;
END bsb

LAYER bsv
  TYPE CUT ;
END bsv

LAYER bm5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 4 ;
  WIDTH 2 ;
  PROPERTY LEF58_WIDTH "WIDTH 2 WRONGDIRECTION ;" ;
END bm5

LAYER bv4
  TYPE CUT ;
END bv4

LAYER bm4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.08 ;
  WIDTH 0.54 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.54 WRONGDIRECTION ;" ;
END bm4

LAYER bv3
  TYPE CUT ;
END bv3

LAYER bm3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.08 ;
  WIDTH 0.54 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.54 WRONGDIRECTION ;" ;
END bm3

LAYER bv2
  TYPE CUT ;
END bv2

LAYER bm2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.38 ;
  WIDTH 0.24 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.24 WRONGDIRECTION ;" ;
END bm2

LAYER bv1
  TYPE CUT ;
END bv1

LAYER bm1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.3 ;
  WIDTH 0.16 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.16 WRONGDIRECTION ;" ;
END bm1

LAYER bv0
  TYPE CUT ;
END bv0

LAYER bm0
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.16 ;
  WIDTH 0.08 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.08 WRONGDIRECTION ;" ;
END bm0

LAYER devflav_n1_id
  TYPE IMPLANT ;
END devflav_n1_id

LAYER vg
  TYPE CUT ;
END vg

LAYER m0
  TYPE ROUTING ;
  MASK 2 ;
  DIRECTION HORIZONTAL ;
  PITCH 0.036 ;
  WIDTH 0.02 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.028 WRONGDIRECTION ;" ;
END m0

LAYER v0
  TYPE CUT ;
END v0

LAYER m1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.05 ;
  WIDTH 0.03 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.035 WRONGDIRECTION ;" ;
END m1

LAYER v1
  TYPE CUT ;
END v1

LAYER m2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.036 ;
  WIDTH 0.02 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END m2

LAYER v2
  TYPE CUT ;
END v2

LAYER m3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.04 ;
  WIDTH 0.024 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END m3

LAYER v3
  TYPE CUT ;
END v3

LAYER m4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.04 ;
  WIDTH 0.024 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END m4

LAYER v4
  TYPE CUT ;
END v4

LAYER m5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.08 ;
  WIDTH 0.04 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.08 WRONGDIRECTION ;" ;
END m5

LAYER v5
  TYPE CUT ;
END v5

LAYER m6
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.08 ;
  WIDTH 0.04 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.08 WRONGDIRECTION ;" ;
END m6

LAYER v6
  TYPE CUT ;
END v6

LAYER m7
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.08 ;
  WIDTH 0.04 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.08 WRONGDIRECTION ;" ;
END m7

LAYER v7
  TYPE CUT ;
END v7

LAYER m8
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.08 ;
  WIDTH 0.04 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.08 WRONGDIRECTION ;" ;
END m8

LAYER v8
  TYPE CUT ;
END v8

LAYER m9
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.08 ;
  WIDTH 0.04 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.08 WRONGDIRECTION ;" ;
END m9

LAYER v9
  TYPE CUT ;
END v9

LAYER m10
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.08 ;
  WIDTH 0.04 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.08 WRONGDIRECTION ;" ;
END m10

LAYER v10
  TYPE CUT ;
END v10

LAYER m11
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.12 ;
  WIDTH 0.06 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.12 WRONGDIRECTION ;" ;
END m11

LAYER v11
  TYPE CUT ;
END v11

LAYER m12
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.12 ;
  WIDTH 0.06 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.12 WRONGDIRECTION ;" ;
END m12

LAYER v12
  TYPE CUT ;
END v12

LAYER m13
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.16 ;
  WIDTH 0.08 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.16 WRONGDIRECTION ;" ;
END m13

LAYER v13
  TYPE CUT ;
END v13

LAYER m14
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.16 ;
  WIDTH 0.08 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.16 WRONGDIRECTION ;" ;
END m14

LAYER ndiff
  TYPE MASTERSLICE ;
END ndiff

LAYER bsbemib
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 45 ;
  WIDTH 20 ;
  PROPERTY LEF58_WIDTH "WIDTH 20 WRONGDIRECTION ;" ;
END bsbemib

LAYER dummy81
  TYPE MASTERSLICE ;
END dummy81

LAYER foundryid
  TYPE MASTERSLICE ;
END foundryid

LAYER bce3
  TYPE MASTERSLICE ;
END bce3

LAYER bce2
  TYPE MASTERSLICE ;
END bce2

LAYER bce1
  TYPE MASTERSLICE ;
END bce1

LAYER dvb
  TYPE MASTERSLICE ;
END dvb

LAYER sdGen
  TYPE MASTERSLICE ;
END sdGen

LAYER pdiff
  TYPE MASTERSLICE ;
END pdiff

LAYER fti
  TYPE MASTERSLICE ;
END fti

LAYER poly
  TYPE MASTERSLICE ;
END poly

LAYER tcn
  TYPE MASTERSLICE ;
END tcn

LAYER vt
  TYPE MASTERSLICE ;
END vt

LAYER gcn
  TYPE MASTERSLICE ;
END gcn

LAYER tfr
  TYPE MASTERSLICE ;
END tfr

LAYER ESD_mask
  TYPE MASTERSLICE ;
END ESD_mask

LAYER NSD_mask
  TYPE MASTERSLICE ;
END NSD_mask

LAYER PSD_mask
  TYPE MASTERSLICE ;
END PSD_mask

LAYER siGen
  TYPE MASTERSLICE ;
END siGen

LAYER bkr
  TYPE MASTERSLICE ;
END bkr

LAYER chkBoundary
  TYPE MASTERSLICE ;
END chkBoundary

LAYER dummy82
  TYPE MASTERSLICE ;
END dummy82

LAYER dummy63
  TYPE MASTERSLICE ;
END dummy63

LAYER dummy273
  TYPE MASTERSLICE ;
END dummy273

LAYER devflav_p1_id
  TYPE IMPLANT ;
END devflav_p1_id

LAYER devflav_n2_id
  TYPE IMPLANT ;
END devflav_n2_id

LAYER devflav_p2_id
  TYPE IMPLANT ;
END devflav_p2_id

LAYER devflav_n3_id
  TYPE IMPLANT ;
END devflav_n3_id

LAYER devflav_p3_id
  TYPE IMPLANT ;
END devflav_p3_id

LAYER devflav_n4_id
  TYPE IMPLANT ;
END devflav_n4_id

LAYER devflav_p4_id
  TYPE IMPLANT ;
END devflav_p4_id

LAYER devflav_n5_id
  TYPE IMPLANT ;
END devflav_n5_id

LAYER devflav_p5_id
  TYPE IMPLANT ;
END devflav_p5_id

VIA BSV_12000x24000_18000V_32000H
  LAYER bsb ;
    RECT -16 -16 16 16 ;
  LAYER bsv ;
    RECT -6 -12 6 12 ;
  LAYER bm5 ;
    RECT -9 -15 9 15 ;
END BSV_12000x24000_18000V_32000H

VIA BSV_12000x24000_18000V_32000V
  LAYER bsb ;
    RECT -16 -16 16 16 ;
  LAYER bsv ;
    RECT -6 -12 6 12 ;
  LAYER bm5 ;
    RECT -9 -15 9 15 ;
END BSV_12000x24000_18000V_32000V

VIA BSV_12000x24000_18000V_35000H
  LAYER bsb ;
    RECT -17.5 -17.5 17.5 17.5 ;
  LAYER bsv ;
    RECT -6 -12 6 12 ;
  LAYER bm5 ;
    RECT -9 -15 9 15 ;
END BSV_12000x24000_18000V_35000H

VIA BSV_12000x24000_18000V_35000V
  LAYER bsb ;
    RECT -17.5 -17.5 17.5 17.5 ;
  LAYER bsv ;
    RECT -6 -12 6 12 ;
  LAYER bm5 ;
    RECT -9 -15 9 15 ;
END BSV_12000x24000_18000V_35000V

VIA BSV_18000x6000_12000H_20000H
  LAYER bsbemib ;
    RECT -10 -10 10 10 ;
  LAYER bsv ;
    RECT -9 -3 9 3 ;
  LAYER bm5 ;
    RECT -12 -6 12 6 ;
END BSV_18000x6000_12000H_20000H

VIA BSV_18000x6000_12000H_20000V
  LAYER bsbemib ;
    RECT -10 -10 10 10 ;
  LAYER bsv ;
    RECT -9 -3 9 3 ;
  LAYER bm5 ;
    RECT -12 -6 12 6 ;
END BSV_18000x6000_12000H_20000V

VIA BSV_18000x6000_24000V_20000H
  LAYER bsbemib ;
    RECT -10 -10 10 10 ;
  LAYER bsv ;
    RECT -9 -3 9 3 ;
  LAYER bm5 ;
    RECT -12 -6 12 6 ;
END BSV_18000x6000_24000V_20000H

VIA BSV_18000x6000_24000V_20000V
  LAYER bsbemib ;
    RECT -10 -10 10 10 ;
  LAYER bsv ;
    RECT -9 -3 9 3 ;
  LAYER bm5 ;
    RECT -12 -6 12 6 ;
END BSV_18000x6000_24000V_20000V

VIA BSV_24000x12000_18000H_32000H
  LAYER bsb ;
    RECT -16 -16 16 16 ;
  LAYER bsv ;
    RECT -12 -6 12 6 ;
  LAYER bm5 ;
    RECT -15 -9 15 9 ;
END BSV_24000x12000_18000H_32000H

VIA BSV_24000x12000_18000H_32000V
  LAYER bsb ;
    RECT -16 -16 16 16 ;
  LAYER bsv ;
    RECT -12 -6 12 6 ;
  LAYER bm5 ;
    RECT -15 -9 15 9 ;
END BSV_24000x12000_18000H_32000V

VIA BSV_24000x12000_18000H_35000H
  LAYER bsb ;
    RECT -17.5 -17.5 17.5 17.5 ;
  LAYER bsv ;
    RECT -12 -6 12 6 ;
  LAYER bm5 ;
    RECT -15 -9 15 9 ;
END BSV_24000x12000_18000H_35000H

VIA BSV_24000x12000_18000H_35000V
  LAYER bsb ;
    RECT -17.5 -17.5 17.5 17.5 ;
  LAYER bsv ;
    RECT -12 -6 12 6 ;
  LAYER bm5 ;
    RECT -15 -9 15 9 ;
END BSV_24000x12000_18000H_35000V

VIA BSV_30000x6000_12000H_51000H
  LAYER bsb ;
    RECT -25.5 -25.5 25.5 25.5 ;
  LAYER bsv ;
    RECT -15 -3 15 3 ;
  LAYER bm5 ;
    RECT -18 -6 18 6 ;
END BSV_30000x6000_12000H_51000H

VIA BSV_30000x6000_12000H_51000V
  LAYER bsb ;
    RECT -25.5 -25.5 25.5 25.5 ;
  LAYER bsv ;
    RECT -15 -3 15 3 ;
  LAYER bm5 ;
    RECT -18 -6 18 6 ;
END BSV_30000x6000_12000H_51000V

VIA BSV_6000x18000_12000V_20000H
  LAYER bsbemib ;
    RECT -10 -10 10 10 ;
  LAYER bsv ;
    RECT -3 -9 3 9 ;
  LAYER bm5 ;
    RECT -6 -12 6 12 ;
END BSV_6000x18000_12000V_20000H

VIA BSV_6000x18000_12000V_20000V
  LAYER bsbemib ;
    RECT -10 -10 10 10 ;
  LAYER bsv ;
    RECT -3 -9 3 9 ;
  LAYER bm5 ;
    RECT -6 -12 6 12 ;
END BSV_6000x18000_12000V_20000V

VIA BSV_6000x18000_24000H_20000H
  LAYER bsbemib ;
    RECT -10 -10 10 10 ;
  LAYER bsv ;
    RECT -3 -9 3 9 ;
  LAYER bm5 ;
    RECT -6 -12 6 12 ;
END BSV_6000x18000_24000H_20000H

VIA BSV_6000x18000_24000H_20000V
  LAYER bsbemib ;
    RECT -10 -10 10 10 ;
  LAYER bsv ;
    RECT -3 -9 3 9 ;
  LAYER bm5 ;
    RECT -6 -12 6 12 ;
END BSV_6000x18000_24000H_20000V

VIA BSV_6000x30000_12000V_51000H
  LAYER bsb ;
    RECT -25.5 -25.5 25.5 25.5 ;
  LAYER bsv ;
    RECT -3 -15 3 15 ;
  LAYER bm5 ;
    RECT -6 -18 6 18 ;
END BSV_6000x30000_12000V_51000H

VIA BSV_6000x30000_12000V_51000V
  LAYER bsb ;
    RECT -25.5 -25.5 25.5 25.5 ;
  LAYER bsv ;
    RECT -3 -15 3 15 ;
  LAYER bm5 ;
    RECT -6 -18 6 18 ;
END BSV_6000x30000_12000V_51000V

VIA BV0_160x260_180V_160V
  LAYER bm1 ;
    RECT -0.08 -0.17 0.08 0.17 ;
  LAYER bv0 ;
    RECT -0.08 -0.13 0.08 0.13 ;
  LAYER bm0 ;
    RECT -0.09 -0.17 0.09 0.17 ;
END BV0_160x260_180V_160V

VIA BV0_160x260_180V_240V
  LAYER bm1 ;
    RECT -0.12 -0.17 0.12 0.17 ;
  LAYER bv0 ;
    RECT -0.08 -0.13 0.08 0.13 ;
  LAYER bm0 ;
    RECT -0.09 -0.17 0.09 0.17 ;
END BV0_160x260_180V_240V

VIA BV0_160x260_180V_320H
  LAYER bm1 ;
    RECT -0.12 -0.16 0.12 0.16 ;
  LAYER bv0 ;
    RECT -0.08 -0.13 0.08 0.13 ;
  LAYER bm0 ;
    RECT -0.09 -0.17 0.09 0.17 ;
END BV0_160x260_180V_320H

VIA BV0_160x260_180V_320V
  LAYER bm1 ;
    RECT -0.16 -0.17 0.16 0.17 ;
  LAYER bv0 ;
    RECT -0.08 -0.13 0.08 0.13 ;
  LAYER bm0 ;
    RECT -0.09 -0.17 0.09 0.17 ;
END BV0_160x260_180V_320V

VIA BV0_160x80_180H_160H
  LAYER bm1 ;
    RECT -0.12 -0.08 0.12 0.08 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END BV0_160x80_180H_160H

VIA BV0_160x80_180H_160V
  LAYER bm1 ;
    RECT -0.08 -0.08 0.08 0.08 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END BV0_160x80_180H_160V

VIA BV0_160x80_180H_240H
  LAYER bm1 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END BV0_160x80_180H_240H

VIA BV0_160x80_180H_240V
  LAYER bm1 ;
    RECT -0.12 -0.08 0.12 0.08 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END BV0_160x80_180H_240V

VIA BV0_160x80_180H_320H
  LAYER bm1 ;
    RECT -0.12 -0.16 0.12 0.16 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END BV0_160x80_180H_320H

VIA BV0_160x80_180H_320V
  LAYER bm1 ;
    RECT -0.16 -0.08 0.16 0.08 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END BV0_160x80_180H_320V

VIA BV0_160x80_180V_160H
  LAYER bm1 ;
    RECT -0.12 -0.08 0.12 0.08 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.09 -0.08 0.09 0.08 ;
END BV0_160x80_180V_160H

VIA BV0_160x80_180V_160V
  LAYER bm1 ;
    RECT -0.08 -0.08 0.08 0.08 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.09 -0.08 0.09 0.08 ;
END BV0_160x80_180V_160V

VIA BV0_160x80_180V_240H
  LAYER bm1 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.09 -0.08 0.09 0.08 ;
END BV0_160x80_180V_240H

VIA BV0_160x80_180V_240V
  LAYER bm1 ;
    RECT -0.12 -0.08 0.12 0.08 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.09 -0.08 0.09 0.08 ;
END BV0_160x80_180V_240V

VIA BV0_160x80_180V_320H
  LAYER bm1 ;
    RECT -0.12 -0.16 0.12 0.16 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.09 -0.08 0.09 0.08 ;
END BV0_160x80_180V_320H

VIA BV0_160x80_180V_320V
  LAYER bm1 ;
    RECT -0.16 -0.08 0.16 0.08 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.09 -0.08 0.09 0.08 ;
END BV0_160x80_180V_320V

VIA BV0_160x80_80H_160H
  LAYER bm1 ;
    RECT -0.12 -0.08 0.12 0.08 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.12 -0.04 0.12 0.04 ;
END BV0_160x80_80H_160H

VIA BV0_160x80_80H_160V
  LAYER bm1 ;
    RECT -0.08 -0.08 0.08 0.08 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.12 -0.04 0.12 0.04 ;
END BV0_160x80_80H_160V

VIA BV0_160x80_80H_240H
  LAYER bm1 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.12 -0.04 0.12 0.04 ;
END BV0_160x80_80H_240H

VIA BV0_160x80_80H_240V
  LAYER bm1 ;
    RECT -0.12 -0.08 0.12 0.08 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.12 -0.04 0.12 0.04 ;
END BV0_160x80_80H_240V

VIA BV0_160x80_80H_320H
  LAYER bm1 ;
    RECT -0.12 -0.16 0.12 0.16 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.12 -0.04 0.12 0.04 ;
END BV0_160x80_80H_320H

VIA BV0_160x80_80H_320V
  LAYER bm1 ;
    RECT -0.16 -0.08 0.16 0.08 ;
  LAYER bv0 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER bm0 ;
    RECT -0.12 -0.04 0.12 0.04 ;
END BV0_160x80_80H_320V

VIA BV0_240x80_180H_160H
  LAYER bm1 ;
    RECT -0.16 -0.08 0.16 0.08 ;
  LAYER bv0 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER bm0 ;
    RECT -0.16 -0.09 0.16 0.09 ;
END BV0_240x80_180H_160H

VIA BV0_240x80_180H_240H
  LAYER bm1 ;
    RECT -0.16 -0.12 0.16 0.12 ;
  LAYER bv0 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER bm0 ;
    RECT -0.16 -0.09 0.16 0.09 ;
END BV0_240x80_180H_240H

VIA BV0_240x80_180H_240V
  LAYER bm1 ;
    RECT -0.12 -0.08 0.12 0.08 ;
  LAYER bv0 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER bm0 ;
    RECT -0.16 -0.09 0.16 0.09 ;
END BV0_240x80_180H_240V

VIA BV0_240x80_180H_320H
  LAYER bm1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER bv0 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER bm0 ;
    RECT -0.16 -0.09 0.16 0.09 ;
END BV0_240x80_180H_320H

VIA BV0_240x80_180H_320V
  LAYER bm1 ;
    RECT -0.16 -0.08 0.16 0.08 ;
  LAYER bv0 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER bm0 ;
    RECT -0.16 -0.09 0.16 0.09 ;
END BV0_240x80_180H_320V

VIA BV0_240x80_80H_160H
  LAYER bm1 ;
    RECT -0.16 -0.08 0.16 0.08 ;
  LAYER bv0 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER bm0 ;
    RECT -0.16 -0.04 0.16 0.04 ;
END BV0_240x80_80H_160H

VIA BV0_240x80_80H_240H
  LAYER bm1 ;
    RECT -0.16 -0.12 0.16 0.12 ;
  LAYER bv0 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER bm0 ;
    RECT -0.16 -0.04 0.16 0.04 ;
END BV0_240x80_80H_240H

VIA BV0_240x80_80H_240V
  LAYER bm1 ;
    RECT -0.12 -0.08 0.12 0.08 ;
  LAYER bv0 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER bm0 ;
    RECT -0.16 -0.04 0.16 0.04 ;
END BV0_240x80_80H_240V

VIA BV0_240x80_80H_320H
  LAYER bm1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER bv0 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER bm0 ;
    RECT -0.16 -0.04 0.16 0.04 ;
END BV0_240x80_80H_320H

VIA BV0_240x80_80H_320V
  LAYER bm1 ;
    RECT -0.16 -0.08 0.16 0.08 ;
  LAYER bv0 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER bm0 ;
    RECT -0.16 -0.04 0.16 0.04 ;
END BV0_240x80_80H_320V

VIA BV0_260x160_180H_160H
  LAYER bm1 ;
    RECT -0.17 -0.08 0.17 0.08 ;
  LAYER bv0 ;
    RECT -0.13 -0.08 0.13 0.08 ;
  LAYER bm0 ;
    RECT -0.17 -0.09 0.17 0.09 ;
END BV0_260x160_180H_160H

VIA BV0_260x160_180H_240H
  LAYER bm1 ;
    RECT -0.17 -0.12 0.17 0.12 ;
  LAYER bv0 ;
    RECT -0.13 -0.08 0.13 0.08 ;
  LAYER bm0 ;
    RECT -0.17 -0.09 0.17 0.09 ;
END BV0_260x160_180H_240H

VIA BV0_260x160_180H_320H
  LAYER bm1 ;
    RECT -0.17 -0.16 0.17 0.16 ;
  LAYER bv0 ;
    RECT -0.13 -0.08 0.13 0.08 ;
  LAYER bm0 ;
    RECT -0.17 -0.09 0.17 0.09 ;
END BV0_260x160_180H_320H

VIA BV0_260x160_180H_320V
  LAYER bm1 ;
    RECT -0.16 -0.12 0.16 0.12 ;
  LAYER bv0 ;
    RECT -0.13 -0.08 0.13 0.08 ;
  LAYER bm0 ;
    RECT -0.17 -0.09 0.17 0.09 ;
END BV0_260x160_180H_320V

VIA BV0_80x160_180H_160H
  LAYER bm1 ;
    RECT -0.08 -0.08 0.08 0.08 ;
  LAYER bv0 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER bm0 ;
    RECT -0.08 -0.09 0.08 0.09 ;
END BV0_80x160_180H_160H

VIA BV0_80x160_180H_160V
  LAYER bm1 ;
    RECT -0.08 -0.12 0.08 0.12 ;
  LAYER bv0 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER bm0 ;
    RECT -0.08 -0.09 0.08 0.09 ;
END BV0_80x160_180H_160V

VIA BV0_80x160_180H_240H
  LAYER bm1 ;
    RECT -0.08 -0.12 0.08 0.12 ;
  LAYER bv0 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER bm0 ;
    RECT -0.08 -0.09 0.08 0.09 ;
END BV0_80x160_180H_240H

VIA BV0_80x160_180H_240V
  LAYER bm1 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER bv0 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER bm0 ;
    RECT -0.08 -0.09 0.08 0.09 ;
END BV0_80x160_180H_240V

VIA BV0_80x160_180H_320H
  LAYER bm1 ;
    RECT -0.08 -0.16 0.08 0.16 ;
  LAYER bv0 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER bm0 ;
    RECT -0.08 -0.09 0.08 0.09 ;
END BV0_80x160_180H_320H

VIA BV0_80x160_180H_320V
  LAYER bm1 ;
    RECT -0.16 -0.12 0.16 0.12 ;
  LAYER bv0 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER bm0 ;
    RECT -0.08 -0.09 0.08 0.09 ;
END BV0_80x160_180H_320V

VIA BV0_80x160_180V_160H
  LAYER bm1 ;
    RECT -0.08 -0.08 0.08 0.08 ;
  LAYER bv0 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER bm0 ;
    RECT -0.09 -0.12 0.09 0.12 ;
END BV0_80x160_180V_160H

VIA BV0_80x160_180V_160V
  LAYER bm1 ;
    RECT -0.08 -0.12 0.08 0.12 ;
  LAYER bv0 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER bm0 ;
    RECT -0.09 -0.12 0.09 0.12 ;
END BV0_80x160_180V_160V

VIA BV0_80x160_180V_240H
  LAYER bm1 ;
    RECT -0.08 -0.12 0.08 0.12 ;
  LAYER bv0 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER bm0 ;
    RECT -0.09 -0.12 0.09 0.12 ;
END BV0_80x160_180V_240H

VIA BV0_80x160_180V_240V
  LAYER bm1 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER bv0 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER bm0 ;
    RECT -0.09 -0.12 0.09 0.12 ;
END BV0_80x160_180V_240V

VIA BV0_80x160_180V_320H
  LAYER bm1 ;
    RECT -0.08 -0.16 0.08 0.16 ;
  LAYER bv0 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER bm0 ;
    RECT -0.09 -0.12 0.09 0.12 ;
END BV0_80x160_180V_320H

VIA BV0_80x160_180V_320V
  LAYER bm1 ;
    RECT -0.16 -0.12 0.16 0.12 ;
  LAYER bv0 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER bm0 ;
    RECT -0.09 -0.12 0.09 0.12 ;
END BV0_80x160_180V_320V

VIA BV0_80x240_180V_160V
  LAYER bm1 ;
    RECT -0.08 -0.16 0.08 0.16 ;
  LAYER bv0 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER bm0 ;
    RECT -0.09 -0.16 0.09 0.16 ;
END BV0_80x240_180V_160V

VIA BV0_80x240_180V_240H
  LAYER bm1 ;
    RECT -0.08 -0.12 0.08 0.12 ;
  LAYER bv0 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER bm0 ;
    RECT -0.09 -0.16 0.09 0.16 ;
END BV0_80x240_180V_240H

VIA BV0_80x240_180V_240V
  LAYER bm1 ;
    RECT -0.12 -0.16 0.12 0.16 ;
  LAYER bv0 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER bm0 ;
    RECT -0.09 -0.16 0.09 0.16 ;
END BV0_80x240_180V_240V

VIA BV0_80x240_180V_320H
  LAYER bm1 ;
    RECT -0.08 -0.16 0.08 0.16 ;
  LAYER bv0 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER bm0 ;
    RECT -0.09 -0.16 0.09 0.16 ;
END BV0_80x240_180V_320H

VIA BV0_80x240_180V_320V
  LAYER bm1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER bv0 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER bm0 ;
    RECT -0.09 -0.16 0.09 0.16 ;
END BV0_80x240_180V_320V

VIA BV1_160x340_160V_240V
  LAYER bm2 ;
    RECT -0.12 -0.29 0.12 0.29 ;
  LAYER bv1 ;
    RECT -0.08 -0.17 0.08 0.17 ;
  LAYER bm1 ;
    RECT -0.08 -0.27 0.08 0.27 ;
END BV1_160x340_160V_240V

VIA BV1_160x340_160V_340H
  LAYER bm2 ;
    RECT -0.2 -0.17 0.2 0.17 ;
  LAYER bv1 ;
    RECT -0.08 -0.17 0.08 0.17 ;
  LAYER bm1 ;
    RECT -0.08 -0.27 0.08 0.27 ;
END BV1_160x340_160V_340H

VIA BV1_160x340_160V_340V
  LAYER bm2 ;
    RECT -0.17 -0.29 0.17 0.29 ;
  LAYER bv1 ;
    RECT -0.08 -0.17 0.08 0.17 ;
  LAYER bm1 ;
    RECT -0.08 -0.27 0.08 0.27 ;
END BV1_160x340_160V_340V

VIA BV1_160x340_160V_510H
  LAYER bm2 ;
    RECT -0.2 -0.255 0.2 0.255 ;
  LAYER bv1 ;
    RECT -0.08 -0.17 0.08 0.17 ;
  LAYER bm1 ;
    RECT -0.08 -0.27 0.08 0.27 ;
END BV1_160x340_160V_510H

VIA BV1_160x340_160V_510V
  LAYER bm2 ;
    RECT -0.255 -0.29 0.255 0.29 ;
  LAYER bv1 ;
    RECT -0.08 -0.17 0.08 0.17 ;
  LAYER bm1 ;
    RECT -0.08 -0.27 0.08 0.27 ;
END BV1_160x340_160V_510V

VIA BV1_160x340_240V_240V
  LAYER bm2 ;
    RECT -0.12 -0.29 0.12 0.29 ;
  LAYER bv1 ;
    RECT -0.08 -0.17 0.08 0.17 ;
  LAYER bm1 ;
    RECT -0.12 -0.27 0.12 0.27 ;
END BV1_160x340_240V_240V

VIA BV1_160x340_240V_340H
  LAYER bm2 ;
    RECT -0.2 -0.17 0.2 0.17 ;
  LAYER bv1 ;
    RECT -0.08 -0.17 0.08 0.17 ;
  LAYER bm1 ;
    RECT -0.12 -0.27 0.12 0.27 ;
END BV1_160x340_240V_340H

VIA BV1_160x340_240V_340V
  LAYER bm2 ;
    RECT -0.17 -0.29 0.17 0.29 ;
  LAYER bv1 ;
    RECT -0.08 -0.17 0.08 0.17 ;
  LAYER bm1 ;
    RECT -0.12 -0.27 0.12 0.27 ;
END BV1_160x340_240V_340V

VIA BV1_160x340_240V_510H
  LAYER bm2 ;
    RECT -0.2 -0.255 0.2 0.255 ;
  LAYER bv1 ;
    RECT -0.08 -0.17 0.08 0.17 ;
  LAYER bm1 ;
    RECT -0.12 -0.27 0.12 0.27 ;
END BV1_160x340_240V_510H

VIA BV1_160x340_240V_510V
  LAYER bm2 ;
    RECT -0.255 -0.29 0.255 0.29 ;
  LAYER bv1 ;
    RECT -0.08 -0.17 0.08 0.17 ;
  LAYER bm1 ;
    RECT -0.12 -0.27 0.12 0.27 ;
END BV1_160x340_240V_510V

VIA BV1_160x340_320V_240V
  LAYER bm2 ;
    RECT -0.12 -0.29 0.12 0.29 ;
  LAYER bv1 ;
    RECT -0.08 -0.17 0.08 0.17 ;
  LAYER bm1 ;
    RECT -0.16 -0.27 0.16 0.27 ;
END BV1_160x340_320V_240V

VIA BV1_160x340_320V_340H
  LAYER bm2 ;
    RECT -0.2 -0.17 0.2 0.17 ;
  LAYER bv1 ;
    RECT -0.08 -0.17 0.08 0.17 ;
  LAYER bm1 ;
    RECT -0.16 -0.27 0.16 0.27 ;
END BV1_160x340_320V_340H

VIA BV1_160x340_320V_340V
  LAYER bm2 ;
    RECT -0.17 -0.29 0.17 0.29 ;
  LAYER bv1 ;
    RECT -0.08 -0.17 0.08 0.17 ;
  LAYER bm1 ;
    RECT -0.16 -0.27 0.16 0.27 ;
END BV1_160x340_320V_340V

VIA BV1_160x340_320V_510H
  LAYER bm2 ;
    RECT -0.2 -0.255 0.2 0.255 ;
  LAYER bv1 ;
    RECT -0.08 -0.17 0.08 0.17 ;
  LAYER bm1 ;
    RECT -0.16 -0.27 0.16 0.27 ;
END BV1_160x340_320V_510H

VIA BV1_160x340_320V_510V
  LAYER bm2 ;
    RECT -0.255 -0.29 0.255 0.29 ;
  LAYER bv1 ;
    RECT -0.08 -0.17 0.08 0.17 ;
  LAYER bm1 ;
    RECT -0.16 -0.27 0.16 0.27 ;
END BV1_160x340_320V_510V

VIA BV1_160x510_160V_240V
  LAYER bm2 ;
    RECT -0.12 -0.375 0.12 0.375 ;
  LAYER bv1 ;
    RECT -0.08 -0.255 0.08 0.255 ;
  LAYER bm1 ;
    RECT -0.08 -0.355 0.08 0.355 ;
END BV1_160x510_160V_240V

VIA BV1_160x510_160V_340V
  LAYER bm2 ;
    RECT -0.17 -0.375 0.17 0.375 ;
  LAYER bv1 ;
    RECT -0.08 -0.255 0.08 0.255 ;
  LAYER bm1 ;
    RECT -0.08 -0.355 0.08 0.355 ;
END BV1_160x510_160V_340V

VIA BV1_160x510_160V_510H
  LAYER bm2 ;
    RECT -0.2 -0.255 0.2 0.255 ;
  LAYER bv1 ;
    RECT -0.08 -0.255 0.08 0.255 ;
  LAYER bm1 ;
    RECT -0.08 -0.355 0.08 0.355 ;
END BV1_160x510_160V_510H

VIA BV1_160x510_160V_510V
  LAYER bm2 ;
    RECT -0.255 -0.375 0.255 0.375 ;
  LAYER bv1 ;
    RECT -0.08 -0.255 0.08 0.255 ;
  LAYER bm1 ;
    RECT -0.08 -0.355 0.08 0.355 ;
END BV1_160x510_160V_510V

VIA BV1_160x510_240V_240V
  LAYER bm2 ;
    RECT -0.12 -0.375 0.12 0.375 ;
  LAYER bv1 ;
    RECT -0.08 -0.255 0.08 0.255 ;
  LAYER bm1 ;
    RECT -0.12 -0.355 0.12 0.355 ;
END BV1_160x510_240V_240V

VIA BV1_160x510_240V_340V
  LAYER bm2 ;
    RECT -0.17 -0.375 0.17 0.375 ;
  LAYER bv1 ;
    RECT -0.08 -0.255 0.08 0.255 ;
  LAYER bm1 ;
    RECT -0.12 -0.355 0.12 0.355 ;
END BV1_160x510_240V_340V

VIA BV1_160x510_240V_510H
  LAYER bm2 ;
    RECT -0.2 -0.255 0.2 0.255 ;
  LAYER bv1 ;
    RECT -0.08 -0.255 0.08 0.255 ;
  LAYER bm1 ;
    RECT -0.12 -0.355 0.12 0.355 ;
END BV1_160x510_240V_510H

VIA BV1_160x510_240V_510V
  LAYER bm2 ;
    RECT -0.255 -0.375 0.255 0.375 ;
  LAYER bv1 ;
    RECT -0.08 -0.255 0.08 0.255 ;
  LAYER bm1 ;
    RECT -0.12 -0.355 0.12 0.355 ;
END BV1_160x510_240V_510V

VIA BV1_160x510_320V_240V
  LAYER bm2 ;
    RECT -0.12 -0.375 0.12 0.375 ;
  LAYER bv1 ;
    RECT -0.08 -0.255 0.08 0.255 ;
  LAYER bm1 ;
    RECT -0.16 -0.355 0.16 0.355 ;
END BV1_160x510_320V_240V

VIA BV1_160x510_320V_340V
  LAYER bm2 ;
    RECT -0.17 -0.375 0.17 0.375 ;
  LAYER bv1 ;
    RECT -0.08 -0.255 0.08 0.255 ;
  LAYER bm1 ;
    RECT -0.16 -0.355 0.16 0.355 ;
END BV1_160x510_320V_340V

VIA BV1_160x510_320V_510H
  LAYER bm2 ;
    RECT -0.2 -0.255 0.2 0.255 ;
  LAYER bv1 ;
    RECT -0.08 -0.255 0.08 0.255 ;
  LAYER bm1 ;
    RECT -0.16 -0.355 0.16 0.355 ;
END BV1_160x510_320V_510H

VIA BV1_160x510_320V_510V
  LAYER bm2 ;
    RECT -0.255 -0.375 0.255 0.375 ;
  LAYER bv1 ;
    RECT -0.08 -0.255 0.08 0.255 ;
  LAYER bm1 ;
    RECT -0.16 -0.355 0.16 0.355 ;
END BV1_160x510_320V_510V

VIA BV1_340x160_160H_240H
  LAYER bm2 ;
    RECT -0.29 -0.12 0.29 0.12 ;
  LAYER bv1 ;
    RECT -0.17 -0.08 0.17 0.08 ;
  LAYER bm1 ;
    RECT -0.27 -0.08 0.27 0.08 ;
END BV1_340x160_160H_240H

VIA BV1_340x160_160H_340H
  LAYER bm2 ;
    RECT -0.29 -0.17 0.29 0.17 ;
  LAYER bv1 ;
    RECT -0.17 -0.08 0.17 0.08 ;
  LAYER bm1 ;
    RECT -0.27 -0.08 0.27 0.08 ;
END BV1_340x160_160H_340H

VIA BV1_340x160_160H_340V
  LAYER bm2 ;
    RECT -0.17 -0.2 0.17 0.2 ;
  LAYER bv1 ;
    RECT -0.17 -0.08 0.17 0.08 ;
  LAYER bm1 ;
    RECT -0.27 -0.08 0.27 0.08 ;
END BV1_340x160_160H_340V

VIA BV1_340x160_160H_510H
  LAYER bm2 ;
    RECT -0.29 -0.255 0.29 0.255 ;
  LAYER bv1 ;
    RECT -0.17 -0.08 0.17 0.08 ;
  LAYER bm1 ;
    RECT -0.27 -0.08 0.27 0.08 ;
END BV1_340x160_160H_510H

VIA BV1_340x160_160H_510V
  LAYER bm2 ;
    RECT -0.255 -0.2 0.255 0.2 ;
  LAYER bv1 ;
    RECT -0.17 -0.08 0.17 0.08 ;
  LAYER bm1 ;
    RECT -0.27 -0.08 0.27 0.08 ;
END BV1_340x160_160H_510V

VIA BV1_340x160_240H_240H
  LAYER bm2 ;
    RECT -0.29 -0.12 0.29 0.12 ;
  LAYER bv1 ;
    RECT -0.17 -0.08 0.17 0.08 ;
  LAYER bm1 ;
    RECT -0.27 -0.12 0.27 0.12 ;
END BV1_340x160_240H_240H

VIA BV1_340x160_240H_340H
  LAYER bm2 ;
    RECT -0.29 -0.17 0.29 0.17 ;
  LAYER bv1 ;
    RECT -0.17 -0.08 0.17 0.08 ;
  LAYER bm1 ;
    RECT -0.27 -0.12 0.27 0.12 ;
END BV1_340x160_240H_340H

VIA BV1_340x160_240H_340V
  LAYER bm2 ;
    RECT -0.17 -0.2 0.17 0.2 ;
  LAYER bv1 ;
    RECT -0.17 -0.08 0.17 0.08 ;
  LAYER bm1 ;
    RECT -0.27 -0.12 0.27 0.12 ;
END BV1_340x160_240H_340V

VIA BV1_340x160_240H_510H
  LAYER bm2 ;
    RECT -0.29 -0.255 0.29 0.255 ;
  LAYER bv1 ;
    RECT -0.17 -0.08 0.17 0.08 ;
  LAYER bm1 ;
    RECT -0.27 -0.12 0.27 0.12 ;
END BV1_340x160_240H_510H

VIA BV1_340x160_240H_510V
  LAYER bm2 ;
    RECT -0.255 -0.2 0.255 0.2 ;
  LAYER bv1 ;
    RECT -0.17 -0.08 0.17 0.08 ;
  LAYER bm1 ;
    RECT -0.27 -0.12 0.27 0.12 ;
END BV1_340x160_240H_510V

VIA BV1_340x160_320H_240H
  LAYER bm2 ;
    RECT -0.29 -0.12 0.29 0.12 ;
  LAYER bv1 ;
    RECT -0.17 -0.08 0.17 0.08 ;
  LAYER bm1 ;
    RECT -0.27 -0.16 0.27 0.16 ;
END BV1_340x160_320H_240H

VIA BV1_340x160_320H_340H
  LAYER bm2 ;
    RECT -0.29 -0.17 0.29 0.17 ;
  LAYER bv1 ;
    RECT -0.17 -0.08 0.17 0.08 ;
  LAYER bm1 ;
    RECT -0.27 -0.16 0.27 0.16 ;
END BV1_340x160_320H_340H

VIA BV1_340x160_320H_340V
  LAYER bm2 ;
    RECT -0.17 -0.2 0.17 0.2 ;
  LAYER bv1 ;
    RECT -0.17 -0.08 0.17 0.08 ;
  LAYER bm1 ;
    RECT -0.27 -0.16 0.27 0.16 ;
END BV1_340x160_320H_340V

VIA BV1_340x160_320H_510H
  LAYER bm2 ;
    RECT -0.29 -0.255 0.29 0.255 ;
  LAYER bv1 ;
    RECT -0.17 -0.08 0.17 0.08 ;
  LAYER bm1 ;
    RECT -0.27 -0.16 0.27 0.16 ;
END BV1_340x160_320H_510H

VIA BV1_340x160_320H_510V
  LAYER bm2 ;
    RECT -0.255 -0.2 0.255 0.2 ;
  LAYER bv1 ;
    RECT -0.17 -0.08 0.17 0.08 ;
  LAYER bm1 ;
    RECT -0.27 -0.16 0.27 0.16 ;
END BV1_340x160_320H_510V

VIA BV1_510x160_160H_240H
  LAYER bm2 ;
    RECT -0.375 -0.12 0.375 0.12 ;
  LAYER bv1 ;
    RECT -0.255 -0.08 0.255 0.08 ;
  LAYER bm1 ;
    RECT -0.355 -0.08 0.355 0.08 ;
END BV1_510x160_160H_240H

VIA BV1_510x160_160H_340H
  LAYER bm2 ;
    RECT -0.375 -0.17 0.375 0.17 ;
  LAYER bv1 ;
    RECT -0.255 -0.08 0.255 0.08 ;
  LAYER bm1 ;
    RECT -0.355 -0.08 0.355 0.08 ;
END BV1_510x160_160H_340H

VIA BV1_510x160_160H_510H
  LAYER bm2 ;
    RECT -0.375 -0.255 0.375 0.255 ;
  LAYER bv1 ;
    RECT -0.255 -0.08 0.255 0.08 ;
  LAYER bm1 ;
    RECT -0.355 -0.08 0.355 0.08 ;
END BV1_510x160_160H_510H

VIA BV1_510x160_160H_510V
  LAYER bm2 ;
    RECT -0.255 -0.2 0.255 0.2 ;
  LAYER bv1 ;
    RECT -0.255 -0.08 0.255 0.08 ;
  LAYER bm1 ;
    RECT -0.355 -0.08 0.355 0.08 ;
END BV1_510x160_160H_510V

VIA BV1_510x160_240H_240H
  LAYER bm2 ;
    RECT -0.375 -0.12 0.375 0.12 ;
  LAYER bv1 ;
    RECT -0.255 -0.08 0.255 0.08 ;
  LAYER bm1 ;
    RECT -0.355 -0.12 0.355 0.12 ;
END BV1_510x160_240H_240H

VIA BV1_510x160_240H_340H
  LAYER bm2 ;
    RECT -0.375 -0.17 0.375 0.17 ;
  LAYER bv1 ;
    RECT -0.255 -0.08 0.255 0.08 ;
  LAYER bm1 ;
    RECT -0.355 -0.12 0.355 0.12 ;
END BV1_510x160_240H_340H

VIA BV1_510x160_240H_510H
  LAYER bm2 ;
    RECT -0.375 -0.255 0.375 0.255 ;
  LAYER bv1 ;
    RECT -0.255 -0.08 0.255 0.08 ;
  LAYER bm1 ;
    RECT -0.355 -0.12 0.355 0.12 ;
END BV1_510x160_240H_510H

VIA BV1_510x160_240H_510V
  LAYER bm2 ;
    RECT -0.255 -0.2 0.255 0.2 ;
  LAYER bv1 ;
    RECT -0.255 -0.08 0.255 0.08 ;
  LAYER bm1 ;
    RECT -0.355 -0.12 0.355 0.12 ;
END BV1_510x160_240H_510V

VIA BV1_510x160_320H_240H
  LAYER bm2 ;
    RECT -0.375 -0.12 0.375 0.12 ;
  LAYER bv1 ;
    RECT -0.255 -0.08 0.255 0.08 ;
  LAYER bm1 ;
    RECT -0.355 -0.16 0.355 0.16 ;
END BV1_510x160_320H_240H

VIA BV1_510x160_320H_340H
  LAYER bm2 ;
    RECT -0.375 -0.17 0.375 0.17 ;
  LAYER bv1 ;
    RECT -0.255 -0.08 0.255 0.08 ;
  LAYER bm1 ;
    RECT -0.355 -0.16 0.355 0.16 ;
END BV1_510x160_320H_340H

VIA BV1_510x160_320H_510H
  LAYER bm2 ;
    RECT -0.375 -0.255 0.375 0.255 ;
  LAYER bv1 ;
    RECT -0.255 -0.08 0.255 0.08 ;
  LAYER bm1 ;
    RECT -0.355 -0.16 0.355 0.16 ;
END BV1_510x160_320H_510H

VIA BV1_510x160_320H_510V
  LAYER bm2 ;
    RECT -0.255 -0.2 0.255 0.2 ;
  LAYER bv1 ;
    RECT -0.255 -0.08 0.255 0.08 ;
  LAYER bm1 ;
    RECT -0.355 -0.16 0.355 0.16 ;
END BV1_510x160_320H_510V

VIA BV2_120x400_340V_540H
  LAYER bm3 ;
    RECT -0.12 -0.27 0.12 0.27 ;
  LAYER bv2 ;
    RECT -0.06 -0.2 0.06 0.2 ;
  LAYER bm2 ;
    RECT -0.17 -0.32 0.17 0.32 ;
END BV2_120x400_340V_540H

VIA BV2_120x400_340V_540V
  LAYER bm3 ;
    RECT -0.27 -0.26 0.27 0.26 ;
  LAYER bv2 ;
    RECT -0.06 -0.2 0.06 0.2 ;
  LAYER bm2 ;
    RECT -0.17 -0.32 0.17 0.32 ;
END BV2_120x400_340V_540V

VIA BV2_120x400_510V_540H
  LAYER bm3 ;
    RECT -0.12 -0.27 0.12 0.27 ;
  LAYER bv2 ;
    RECT -0.06 -0.2 0.06 0.2 ;
  LAYER bm2 ;
    RECT -0.255 -0.32 0.255 0.32 ;
END BV2_120x400_510V_540H

VIA BV2_120x400_510V_540V
  LAYER bm3 ;
    RECT -0.27 -0.26 0.27 0.26 ;
  LAYER bv2 ;
    RECT -0.06 -0.2 0.06 0.2 ;
  LAYER bm2 ;
    RECT -0.255 -0.32 0.255 0.32 ;
END BV2_120x400_510V_540V

VIA BV2_200x640_340V_540V
  LAYER bm3 ;
    RECT -0.27 -0.38 0.27 0.38 ;
  LAYER bv2 ;
    RECT -0.1 -0.32 0.1 0.32 ;
  LAYER bm2 ;
    RECT -0.17 -0.38 0.17 0.38 ;
END BV2_200x640_340V_540V

VIA BV2_200x640_340V_748H
  LAYER bm3 ;
    RECT -0.16 -0.374 0.16 0.374 ;
  LAYER bv2 ;
    RECT -0.1 -0.32 0.1 0.32 ;
  LAYER bm2 ;
    RECT -0.17 -0.38 0.17 0.38 ;
END BV2_200x640_340V_748H

VIA BV2_200x640_510V_540V
  LAYER bm3 ;
    RECT -0.27 -0.38 0.27 0.38 ;
  LAYER bv2 ;
    RECT -0.1 -0.32 0.1 0.32 ;
  LAYER bm2 ;
    RECT -0.255 -0.38 0.255 0.38 ;
END BV2_200x640_510V_540V

VIA BV2_200x640_510V_748H
  LAYER bm3 ;
    RECT -0.16 -0.374 0.16 0.374 ;
  LAYER bv2 ;
    RECT -0.1 -0.32 0.1 0.32 ;
  LAYER bm2 ;
    RECT -0.255 -0.38 0.255 0.38 ;
END BV2_200x640_510V_748H

VIA BV2_400x120_340H_540H
  LAYER bm3 ;
    RECT -0.26 -0.27 0.26 0.27 ;
  LAYER bv2 ;
    RECT -0.2 -0.06 0.2 0.06 ;
  LAYER bm2 ;
    RECT -0.32 -0.17 0.32 0.17 ;
END BV2_400x120_340H_540H

VIA BV2_400x120_340H_540V
  LAYER bm3 ;
    RECT -0.27 -0.12 0.27 0.12 ;
  LAYER bv2 ;
    RECT -0.2 -0.06 0.2 0.06 ;
  LAYER bm2 ;
    RECT -0.32 -0.17 0.32 0.17 ;
END BV2_400x120_340H_540V

VIA BV2_400x120_510H_540H
  LAYER bm3 ;
    RECT -0.26 -0.27 0.26 0.27 ;
  LAYER bv2 ;
    RECT -0.2 -0.06 0.2 0.06 ;
  LAYER bm2 ;
    RECT -0.32 -0.255 0.32 0.255 ;
END BV2_400x120_510H_540H

VIA BV2_400x120_510H_540V
  LAYER bm3 ;
    RECT -0.27 -0.12 0.27 0.12 ;
  LAYER bv2 ;
    RECT -0.2 -0.06 0.2 0.06 ;
  LAYER bm2 ;
    RECT -0.32 -0.255 0.32 0.255 ;
END BV2_400x120_510H_540V

VIA BV2_640x200_340H_540H
  LAYER bm3 ;
    RECT -0.38 -0.27 0.38 0.27 ;
  LAYER bv2 ;
    RECT -0.32 -0.1 0.32 0.1 ;
  LAYER bm2 ;
    RECT -0.38 -0.17 0.38 0.17 ;
END BV2_640x200_340H_540H

VIA BV2_640x200_340H_748V
  LAYER bm3 ;
    RECT -0.374 -0.16 0.374 0.16 ;
  LAYER bv2 ;
    RECT -0.32 -0.1 0.32 0.1 ;
  LAYER bm2 ;
    RECT -0.38 -0.17 0.38 0.17 ;
END BV2_640x200_340H_748V

VIA BV2_640x200_510H_540H
  LAYER bm3 ;
    RECT -0.38 -0.27 0.38 0.27 ;
  LAYER bv2 ;
    RECT -0.32 -0.1 0.32 0.1 ;
  LAYER bm2 ;
    RECT -0.38 -0.255 0.38 0.255 ;
END BV2_640x200_510H_540H

VIA BV2_640x200_510H_748V
  LAYER bm3 ;
    RECT -0.374 -0.16 0.374 0.16 ;
  LAYER bv2 ;
    RECT -0.32 -0.1 0.32 0.1 ;
  LAYER bm2 ;
    RECT -0.38 -0.255 0.38 0.255 ;
END BV2_640x200_510H_748V

VIA BV3_1200x400_1400V_1200d5H
  LAYER bm4 ;
    RECT -0.72 -0.6 0.72 0.6 ;
  LAYER bv3 ;
    RECT -0.6 -0.2 0.6 0.2 ;
  LAYER bm3 ;
    RECT -0.7 -0.3 0.7 0.3 ;
END BV3_1200x400_1400V_1200d5H

VIA BV3_1200x400_1400V_1440V
  LAYER bm4 ;
    RECT -0.72 -0.32 0.72 0.32 ;
  LAYER bv3 ;
    RECT -0.6 -0.2 0.6 0.2 ;
  LAYER bm3 ;
    RECT -0.7 -0.3 0.7 0.3 ;
END BV3_1200x400_1400V_1440V

VIA BV3_1200x400_1400V_2400d5H
  LAYER bm4 ;
    RECT -0.77 -1.2 0.77 1.2 ;
  LAYER bv3 ;
    RECT -0.6 -0.2 0.6 0.2 ;
  LAYER bm3 ;
    RECT -0.7 -0.3 0.7 0.3 ;
END BV3_1200x400_1400V_2400d5H

VIA BV3_1200x400_1400V_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.37 1.2 0.37 ;
  LAYER bv3 ;
    RECT -0.6 -0.2 0.6 0.2 ;
  LAYER bm3 ;
    RECT -0.7 -0.3 0.7 0.3 ;
END BV3_1200x400_1400V_2400d5V

VIA BV3_1200x400_1400V_540H
  LAYER bm4 ;
    RECT -0.66 -0.27 0.66 0.27 ;
  LAYER bv3 ;
    RECT -0.6 -0.2 0.6 0.2 ;
  LAYER bm3 ;
    RECT -0.7 -0.3 0.7 0.3 ;
END BV3_1200x400_1400V_540H

VIA BV3_1200x400_1400V_720d5H
  LAYER bm4 ;
    RECT -0.685 -0.36 0.685 0.36 ;
  LAYER bv3 ;
    RECT -0.6 -0.2 0.6 0.2 ;
  LAYER bm3 ;
    RECT -0.7 -0.3 0.7 0.3 ;
END BV3_1200x400_1400V_720d5H

VIA BV3_1200x400_600H_1200d5H
  LAYER bm4 ;
    RECT -0.72 -0.6 0.72 0.6 ;
  LAYER bv3 ;
    RECT -0.6 -0.2 0.6 0.2 ;
  LAYER bm3 ;
    RECT -0.7 -0.3 0.7 0.3 ;
END BV3_1200x400_600H_1200d5H

VIA BV3_1200x400_600H_1440V
  LAYER bm4 ;
    RECT -0.72 -0.32 0.72 0.32 ;
  LAYER bv3 ;
    RECT -0.6 -0.2 0.6 0.2 ;
  LAYER bm3 ;
    RECT -0.7 -0.3 0.7 0.3 ;
END BV3_1200x400_600H_1440V

VIA BV3_1200x400_600H_2400d5H
  LAYER bm4 ;
    RECT -0.77 -1.2 0.77 1.2 ;
  LAYER bv3 ;
    RECT -0.6 -0.2 0.6 0.2 ;
  LAYER bm3 ;
    RECT -0.7 -0.3 0.7 0.3 ;
END BV3_1200x400_600H_2400d5H

VIA BV3_1200x400_600H_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.37 1.2 0.37 ;
  LAYER bv3 ;
    RECT -0.6 -0.2 0.6 0.2 ;
  LAYER bm3 ;
    RECT -0.7 -0.3 0.7 0.3 ;
END BV3_1200x400_600H_2400d5V

VIA BV3_1200x400_600H_540H
  LAYER bm4 ;
    RECT -0.66 -0.27 0.66 0.27 ;
  LAYER bv3 ;
    RECT -0.6 -0.2 0.6 0.2 ;
  LAYER bm3 ;
    RECT -0.7 -0.3 0.7 0.3 ;
END BV3_1200x400_600H_540H

VIA BV3_1200x400_600H_720d5H
  LAYER bm4 ;
    RECT -0.685 -0.36 0.685 0.36 ;
  LAYER bv3 ;
    RECT -0.6 -0.2 0.6 0.2 ;
  LAYER bm3 ;
    RECT -0.7 -0.3 0.7 0.3 ;
END BV3_1200x400_600H_720d5H

VIA BV3_1500x400_1700V_1200d5H
  LAYER bm4 ;
    RECT -0.87 -0.6 0.87 0.6 ;
  LAYER bv3 ;
    RECT -0.75 -0.2 0.75 0.2 ;
  LAYER bm3 ;
    RECT -0.85 -0.3 0.85 0.3 ;
END BV3_1500x400_1700V_1200d5H

VIA BV3_1500x400_1700V_1740V
  LAYER bm4 ;
    RECT -0.87 -0.32 0.87 0.32 ;
  LAYER bv3 ;
    RECT -0.75 -0.2 0.75 0.2 ;
  LAYER bm3 ;
    RECT -0.85 -0.3 0.85 0.3 ;
END BV3_1500x400_1700V_1740V

VIA BV3_1500x400_1700V_2400d5H
  LAYER bm4 ;
    RECT -0.92 -1.2 0.92 1.2 ;
  LAYER bv3 ;
    RECT -0.75 -0.2 0.75 0.2 ;
  LAYER bm3 ;
    RECT -0.85 -0.3 0.85 0.3 ;
END BV3_1500x400_1700V_2400d5H

VIA BV3_1500x400_1700V_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.37 1.2 0.37 ;
  LAYER bv3 ;
    RECT -0.75 -0.2 0.75 0.2 ;
  LAYER bm3 ;
    RECT -0.85 -0.3 0.85 0.3 ;
END BV3_1500x400_1700V_2400d5V

VIA BV3_1500x400_1700V_540H
  LAYER bm4 ;
    RECT -0.81 -0.27 0.81 0.27 ;
  LAYER bv3 ;
    RECT -0.75 -0.2 0.75 0.2 ;
  LAYER bm3 ;
    RECT -0.85 -0.3 0.85 0.3 ;
END BV3_1500x400_1700V_540H

VIA BV3_1500x400_1700V_720d5H
  LAYER bm4 ;
    RECT -0.835 -0.36 0.835 0.36 ;
  LAYER bv3 ;
    RECT -0.75 -0.2 0.75 0.2 ;
  LAYER bm3 ;
    RECT -0.85 -0.3 0.85 0.3 ;
END BV3_1500x400_1700V_720d5H

VIA BV3_1500x400_600H_1200d5H
  LAYER bm4 ;
    RECT -0.87 -0.6 0.87 0.6 ;
  LAYER bv3 ;
    RECT -0.75 -0.2 0.75 0.2 ;
  LAYER bm3 ;
    RECT -0.85 -0.3 0.85 0.3 ;
END BV3_1500x400_600H_1200d5H

VIA BV3_1500x400_600H_1740V
  LAYER bm4 ;
    RECT -0.87 -0.32 0.87 0.32 ;
  LAYER bv3 ;
    RECT -0.75 -0.2 0.75 0.2 ;
  LAYER bm3 ;
    RECT -0.85 -0.3 0.85 0.3 ;
END BV3_1500x400_600H_1740V

VIA BV3_1500x400_600H_2400d5H
  LAYER bm4 ;
    RECT -0.92 -1.2 0.92 1.2 ;
  LAYER bv3 ;
    RECT -0.75 -0.2 0.75 0.2 ;
  LAYER bm3 ;
    RECT -0.85 -0.3 0.85 0.3 ;
END BV3_1500x400_600H_2400d5H

VIA BV3_1500x400_600H_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.37 1.2 0.37 ;
  LAYER bv3 ;
    RECT -0.75 -0.2 0.75 0.2 ;
  LAYER bm3 ;
    RECT -0.85 -0.3 0.85 0.3 ;
END BV3_1500x400_600H_2400d5V

VIA BV3_1500x400_600H_540H
  LAYER bm4 ;
    RECT -0.81 -0.27 0.81 0.27 ;
  LAYER bv3 ;
    RECT -0.75 -0.2 0.75 0.2 ;
  LAYER bm3 ;
    RECT -0.85 -0.3 0.85 0.3 ;
END BV3_1500x400_600H_540H

VIA BV3_1500x400_600H_720d5H
  LAYER bm4 ;
    RECT -0.835 -0.36 0.835 0.36 ;
  LAYER bv3 ;
    RECT -0.75 -0.2 0.75 0.2 ;
  LAYER bm3 ;
    RECT -0.85 -0.3 0.85 0.3 ;
END BV3_1500x400_600H_720d5H

VIA BV3_3000x400_3200V_1200d5H
  LAYER bm4 ;
    RECT -1.62 -0.6 1.62 0.6 ;
  LAYER bv3 ;
    RECT -1.5 -0.2 1.5 0.2 ;
  LAYER bm3 ;
    RECT -1.6 -0.3 1.6 0.3 ;
END BV3_3000x400_3200V_1200d5H

VIA BV3_3000x400_3200V_2400d5H
  LAYER bm4 ;
    RECT -1.67 -1.2 1.67 1.2 ;
  LAYER bv3 ;
    RECT -1.5 -0.2 1.5 0.2 ;
  LAYER bm3 ;
    RECT -1.6 -0.3 1.6 0.3 ;
END BV3_3000x400_3200V_2400d5H

VIA BV3_3000x400_3200V_3340V
  LAYER bm4 ;
    RECT -1.67 -0.37 1.67 0.37 ;
  LAYER bv3 ;
    RECT -1.5 -0.2 1.5 0.2 ;
  LAYER bm3 ;
    RECT -1.6 -0.3 1.6 0.3 ;
END BV3_3000x400_3200V_3340V

VIA BV3_3000x400_3200V_540H
  LAYER bm4 ;
    RECT -1.56 -0.27 1.56 0.27 ;
  LAYER bv3 ;
    RECT -1.5 -0.2 1.5 0.2 ;
  LAYER bm3 ;
    RECT -1.6 -0.3 1.6 0.3 ;
END BV3_3000x400_3200V_540H

VIA BV3_3000x400_3200V_720d5H
  LAYER bm4 ;
    RECT -1.585 -0.36 1.585 0.36 ;
  LAYER bv3 ;
    RECT -1.5 -0.2 1.5 0.2 ;
  LAYER bm3 ;
    RECT -1.6 -0.3 1.6 0.3 ;
END BV3_3000x400_3200V_720d5H

VIA BV3_3000x400_600H_1200d5H
  LAYER bm4 ;
    RECT -1.62 -0.6 1.62 0.6 ;
  LAYER bv3 ;
    RECT -1.5 -0.2 1.5 0.2 ;
  LAYER bm3 ;
    RECT -1.6 -0.3 1.6 0.3 ;
END BV3_3000x400_600H_1200d5H

VIA BV3_3000x400_600H_2400d5H
  LAYER bm4 ;
    RECT -1.67 -1.2 1.67 1.2 ;
  LAYER bv3 ;
    RECT -1.5 -0.2 1.5 0.2 ;
  LAYER bm3 ;
    RECT -1.6 -0.3 1.6 0.3 ;
END BV3_3000x400_600H_2400d5H

VIA BV3_3000x400_600H_3340V
  LAYER bm4 ;
    RECT -1.67 -0.37 1.67 0.37 ;
  LAYER bv3 ;
    RECT -1.5 -0.2 1.5 0.2 ;
  LAYER bm3 ;
    RECT -1.6 -0.3 1.6 0.3 ;
END BV3_3000x400_600H_3340V

VIA BV3_3000x400_600H_540H
  LAYER bm4 ;
    RECT -1.56 -0.27 1.56 0.27 ;
  LAYER bv3 ;
    RECT -1.5 -0.2 1.5 0.2 ;
  LAYER bm3 ;
    RECT -1.6 -0.3 1.6 0.3 ;
END BV3_3000x400_600H_540H

VIA BV3_3000x400_600H_720d5H
  LAYER bm4 ;
    RECT -1.585 -0.36 1.585 0.36 ;
  LAYER bv3 ;
    RECT -1.5 -0.2 1.5 0.2 ;
  LAYER bm3 ;
    RECT -1.6 -0.3 1.6 0.3 ;
END BV3_3000x400_600H_720d5H

VIA BV3_400x1200_1400H_1200d5V
  LAYER bm4 ;
    RECT -0.6 -0.72 0.6 0.72 ;
  LAYER bv3 ;
    RECT -0.2 -0.6 0.2 0.6 ;
  LAYER bm3 ;
    RECT -0.3 -0.7 0.3 0.7 ;
END BV3_400x1200_1400H_1200d5V

VIA BV3_400x1200_1400H_1440H
  LAYER bm4 ;
    RECT -0.32 -0.72 0.32 0.72 ;
  LAYER bv3 ;
    RECT -0.2 -0.6 0.2 0.6 ;
  LAYER bm3 ;
    RECT -0.3 -0.7 0.3 0.7 ;
END BV3_400x1200_1400H_1440H

VIA BV3_400x1200_1400H_2400d5H
  LAYER bm4 ;
    RECT -0.37 -1.2 0.37 1.2 ;
  LAYER bv3 ;
    RECT -0.2 -0.6 0.2 0.6 ;
  LAYER bm3 ;
    RECT -0.3 -0.7 0.3 0.7 ;
END BV3_400x1200_1400H_2400d5H

VIA BV3_400x1200_1400H_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.77 1.2 0.77 ;
  LAYER bv3 ;
    RECT -0.2 -0.6 0.2 0.6 ;
  LAYER bm3 ;
    RECT -0.3 -0.7 0.3 0.7 ;
END BV3_400x1200_1400H_2400d5V

VIA BV3_400x1200_1400H_540V
  LAYER bm4 ;
    RECT -0.27 -0.66 0.27 0.66 ;
  LAYER bv3 ;
    RECT -0.2 -0.6 0.2 0.6 ;
  LAYER bm3 ;
    RECT -0.3 -0.7 0.3 0.7 ;
END BV3_400x1200_1400H_540V

VIA BV3_400x1200_1400H_720d5V
  LAYER bm4 ;
    RECT -0.36 -0.685 0.36 0.685 ;
  LAYER bv3 ;
    RECT -0.2 -0.6 0.2 0.6 ;
  LAYER bm3 ;
    RECT -0.3 -0.7 0.3 0.7 ;
END BV3_400x1200_1400H_720d5V

VIA BV3_400x1200_600V_1200d5V
  LAYER bm4 ;
    RECT -0.6 -0.72 0.6 0.72 ;
  LAYER bv3 ;
    RECT -0.2 -0.6 0.2 0.6 ;
  LAYER bm3 ;
    RECT -0.3 -0.7 0.3 0.7 ;
END BV3_400x1200_600V_1200d5V

VIA BV3_400x1200_600V_1440H
  LAYER bm4 ;
    RECT -0.32 -0.72 0.32 0.72 ;
  LAYER bv3 ;
    RECT -0.2 -0.6 0.2 0.6 ;
  LAYER bm3 ;
    RECT -0.3 -0.7 0.3 0.7 ;
END BV3_400x1200_600V_1440H

VIA BV3_400x1200_600V_2400d5H
  LAYER bm4 ;
    RECT -0.37 -1.2 0.37 1.2 ;
  LAYER bv3 ;
    RECT -0.2 -0.6 0.2 0.6 ;
  LAYER bm3 ;
    RECT -0.3 -0.7 0.3 0.7 ;
END BV3_400x1200_600V_2400d5H

VIA BV3_400x1200_600V_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.77 1.2 0.77 ;
  LAYER bv3 ;
    RECT -0.2 -0.6 0.2 0.6 ;
  LAYER bm3 ;
    RECT -0.3 -0.7 0.3 0.7 ;
END BV3_400x1200_600V_2400d5V

VIA BV3_400x1200_600V_540V
  LAYER bm4 ;
    RECT -0.27 -0.66 0.27 0.66 ;
  LAYER bv3 ;
    RECT -0.2 -0.6 0.2 0.6 ;
  LAYER bm3 ;
    RECT -0.3 -0.7 0.3 0.7 ;
END BV3_400x1200_600V_540V

VIA BV3_400x1200_600V_720d5V
  LAYER bm4 ;
    RECT -0.36 -0.685 0.36 0.685 ;
  LAYER bv3 ;
    RECT -0.2 -0.6 0.2 0.6 ;
  LAYER bm3 ;
    RECT -0.3 -0.7 0.3 0.7 ;
END BV3_400x1200_600V_720d5V

VIA BV3_400x1500_1700H_1200d5V
  LAYER bm4 ;
    RECT -0.6 -0.87 0.6 0.87 ;
  LAYER bv3 ;
    RECT -0.2 -0.75 0.2 0.75 ;
  LAYER bm3 ;
    RECT -0.3 -0.85 0.3 0.85 ;
END BV3_400x1500_1700H_1200d5V

VIA BV3_400x1500_1700H_1740H
  LAYER bm4 ;
    RECT -0.32 -0.87 0.32 0.87 ;
  LAYER bv3 ;
    RECT -0.2 -0.75 0.2 0.75 ;
  LAYER bm3 ;
    RECT -0.3 -0.85 0.3 0.85 ;
END BV3_400x1500_1700H_1740H

VIA BV3_400x1500_1700H_2400d5H
  LAYER bm4 ;
    RECT -0.37 -1.2 0.37 1.2 ;
  LAYER bv3 ;
    RECT -0.2 -0.75 0.2 0.75 ;
  LAYER bm3 ;
    RECT -0.3 -0.85 0.3 0.85 ;
END BV3_400x1500_1700H_2400d5H

VIA BV3_400x1500_1700H_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.92 1.2 0.92 ;
  LAYER bv3 ;
    RECT -0.2 -0.75 0.2 0.75 ;
  LAYER bm3 ;
    RECT -0.3 -0.85 0.3 0.85 ;
END BV3_400x1500_1700H_2400d5V

VIA BV3_400x1500_1700H_540V
  LAYER bm4 ;
    RECT -0.27 -0.81 0.27 0.81 ;
  LAYER bv3 ;
    RECT -0.2 -0.75 0.2 0.75 ;
  LAYER bm3 ;
    RECT -0.3 -0.85 0.3 0.85 ;
END BV3_400x1500_1700H_540V

VIA BV3_400x1500_1700H_720d5V
  LAYER bm4 ;
    RECT -0.36 -0.835 0.36 0.835 ;
  LAYER bv3 ;
    RECT -0.2 -0.75 0.2 0.75 ;
  LAYER bm3 ;
    RECT -0.3 -0.85 0.3 0.85 ;
END BV3_400x1500_1700H_720d5V

VIA BV3_400x1500_600V_1200d5V
  LAYER bm4 ;
    RECT -0.6 -0.87 0.6 0.87 ;
  LAYER bv3 ;
    RECT -0.2 -0.75 0.2 0.75 ;
  LAYER bm3 ;
    RECT -0.3 -0.85 0.3 0.85 ;
END BV3_400x1500_600V_1200d5V

VIA BV3_400x1500_600V_1740H
  LAYER bm4 ;
    RECT -0.32 -0.87 0.32 0.87 ;
  LAYER bv3 ;
    RECT -0.2 -0.75 0.2 0.75 ;
  LAYER bm3 ;
    RECT -0.3 -0.85 0.3 0.85 ;
END BV3_400x1500_600V_1740H

VIA BV3_400x1500_600V_2400d5H
  LAYER bm4 ;
    RECT -0.37 -1.2 0.37 1.2 ;
  LAYER bv3 ;
    RECT -0.2 -0.75 0.2 0.75 ;
  LAYER bm3 ;
    RECT -0.3 -0.85 0.3 0.85 ;
END BV3_400x1500_600V_2400d5H

VIA BV3_400x1500_600V_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.92 1.2 0.92 ;
  LAYER bv3 ;
    RECT -0.2 -0.75 0.2 0.75 ;
  LAYER bm3 ;
    RECT -0.3 -0.85 0.3 0.85 ;
END BV3_400x1500_600V_2400d5V

VIA BV3_400x1500_600V_540V
  LAYER bm4 ;
    RECT -0.27 -0.81 0.27 0.81 ;
  LAYER bv3 ;
    RECT -0.2 -0.75 0.2 0.75 ;
  LAYER bm3 ;
    RECT -0.3 -0.85 0.3 0.85 ;
END BV3_400x1500_600V_540V

VIA BV3_400x1500_600V_720d5V
  LAYER bm4 ;
    RECT -0.36 -0.835 0.36 0.835 ;
  LAYER bv3 ;
    RECT -0.2 -0.75 0.2 0.75 ;
  LAYER bm3 ;
    RECT -0.3 -0.85 0.3 0.85 ;
END BV3_400x1500_600V_720d5V

VIA BV3_400x3000_3200H_1200d5V
  LAYER bm4 ;
    RECT -0.6 -1.62 0.6 1.62 ;
  LAYER bv3 ;
    RECT -0.2 -1.5 0.2 1.5 ;
  LAYER bm3 ;
    RECT -0.3 -1.6 0.3 1.6 ;
END BV3_400x3000_3200H_1200d5V

VIA BV3_400x3000_3200H_2400d5V
  LAYER bm4 ;
    RECT -1.2 -1.67 1.2 1.67 ;
  LAYER bv3 ;
    RECT -0.2 -1.5 0.2 1.5 ;
  LAYER bm3 ;
    RECT -0.3 -1.6 0.3 1.6 ;
END BV3_400x3000_3200H_2400d5V

VIA BV3_400x3000_3200H_3340H
  LAYER bm4 ;
    RECT -0.37 -1.67 0.37 1.67 ;
  LAYER bv3 ;
    RECT -0.2 -1.5 0.2 1.5 ;
  LAYER bm3 ;
    RECT -0.3 -1.6 0.3 1.6 ;
END BV3_400x3000_3200H_3340H

VIA BV3_400x3000_3200H_540V
  LAYER bm4 ;
    RECT -0.27 -1.56 0.27 1.56 ;
  LAYER bv3 ;
    RECT -0.2 -1.5 0.2 1.5 ;
  LAYER bm3 ;
    RECT -0.3 -1.6 0.3 1.6 ;
END BV3_400x3000_3200H_540V

VIA BV3_400x3000_3200H_720d5V
  LAYER bm4 ;
    RECT -0.36 -1.585 0.36 1.585 ;
  LAYER bv3 ;
    RECT -0.2 -1.5 0.2 1.5 ;
  LAYER bm3 ;
    RECT -0.3 -1.6 0.3 1.6 ;
END BV3_400x3000_3200H_720d5V

VIA BV3_400x3000_600V_1200d5V
  LAYER bm4 ;
    RECT -0.6 -1.62 0.6 1.62 ;
  LAYER bv3 ;
    RECT -0.2 -1.5 0.2 1.5 ;
  LAYER bm3 ;
    RECT -0.3 -1.6 0.3 1.6 ;
END BV3_400x3000_600V_1200d5V

VIA BV3_400x3000_600V_2400d5V
  LAYER bm4 ;
    RECT -1.2 -1.67 1.2 1.67 ;
  LAYER bv3 ;
    RECT -0.2 -1.5 0.2 1.5 ;
  LAYER bm3 ;
    RECT -0.3 -1.6 0.3 1.6 ;
END BV3_400x3000_600V_2400d5V

VIA BV3_400x3000_600V_3340H
  LAYER bm4 ;
    RECT -0.37 -1.67 0.37 1.67 ;
  LAYER bv3 ;
    RECT -0.2 -1.5 0.2 1.5 ;
  LAYER bm3 ;
    RECT -0.3 -1.6 0.3 1.6 ;
END BV3_400x3000_600V_3340H

VIA BV3_400x3000_600V_540V
  LAYER bm4 ;
    RECT -0.27 -1.56 0.27 1.56 ;
  LAYER bv3 ;
    RECT -0.2 -1.5 0.2 1.5 ;
  LAYER bm3 ;
    RECT -0.3 -1.6 0.3 1.6 ;
END BV3_400x3000_600V_540V

VIA BV3_400x3000_600V_720d5V
  LAYER bm4 ;
    RECT -0.36 -1.585 0.36 1.585 ;
  LAYER bv3 ;
    RECT -0.2 -1.5 0.2 1.5 ;
  LAYER bm3 ;
    RECT -0.3 -1.6 0.3 1.6 ;
END BV3_400x3000_600V_720d5V

VIA BV3_400x400_540H_1200d5H
  LAYER bm4 ;
    RECT -0.32 -0.6 0.32 0.6 ;
  LAYER bv3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER bm3 ;
    RECT -0.27 -0.27 0.27 0.27 ;
END BV3_400x400_540H_1200d5H

VIA BV3_400x400_540H_1200d5V
  LAYER bm4 ;
    RECT -0.6 -0.32 0.6 0.32 ;
  LAYER bv3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER bm3 ;
    RECT -0.27 -0.27 0.27 0.27 ;
END BV3_400x400_540H_1200d5V

VIA BV3_400x400_540H_2400d5H
  LAYER bm4 ;
    RECT -0.37 -1.2 0.37 1.2 ;
  LAYER bv3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER bm3 ;
    RECT -0.27 -0.27 0.27 0.27 ;
END BV3_400x400_540H_2400d5H

VIA BV3_400x400_540H_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.37 1.2 0.37 ;
  LAYER bv3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER bm3 ;
    RECT -0.27 -0.27 0.27 0.27 ;
END BV3_400x400_540H_2400d5V

VIA BV3_400x400_540H_540H
  LAYER bm4 ;
    RECT -0.26 -0.27 0.26 0.27 ;
  LAYER bv3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER bm3 ;
    RECT -0.27 -0.27 0.27 0.27 ;
END BV3_400x400_540H_540H

VIA BV3_400x400_540H_540V
  LAYER bm4 ;
    RECT -0.27 -0.26 0.27 0.26 ;
  LAYER bv3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER bm3 ;
    RECT -0.27 -0.27 0.27 0.27 ;
END BV3_400x400_540H_540V

VIA BV3_400x400_540H_720d5H
  LAYER bm4 ;
    RECT -0.285 -0.36 0.285 0.36 ;
  LAYER bv3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER bm3 ;
    RECT -0.27 -0.27 0.27 0.27 ;
END BV3_400x400_540H_720d5H

VIA BV3_400x400_540H_720d5V
  LAYER bm4 ;
    RECT -0.36 -0.285 0.36 0.285 ;
  LAYER bv3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER bm3 ;
    RECT -0.27 -0.27 0.27 0.27 ;
END BV3_400x400_540H_720d5V

VIA BV3_400x400_540V_1200d5H
  LAYER bm4 ;
    RECT -0.32 -0.6 0.32 0.6 ;
  LAYER bv3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER bm3 ;
    RECT -0.27 -0.27 0.27 0.27 ;
END BV3_400x400_540V_1200d5H

VIA BV3_400x400_540V_1200d5V
  LAYER bm4 ;
    RECT -0.6 -0.32 0.6 0.32 ;
  LAYER bv3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER bm3 ;
    RECT -0.27 -0.27 0.27 0.27 ;
END BV3_400x400_540V_1200d5V

VIA BV3_400x400_540V_2400d5H
  LAYER bm4 ;
    RECT -0.37 -1.2 0.37 1.2 ;
  LAYER bv3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER bm3 ;
    RECT -0.27 -0.27 0.27 0.27 ;
END BV3_400x400_540V_2400d5H

VIA BV3_400x400_540V_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.37 1.2 0.37 ;
  LAYER bv3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER bm3 ;
    RECT -0.27 -0.27 0.27 0.27 ;
END BV3_400x400_540V_2400d5V

VIA BV3_400x400_540V_540H
  LAYER bm4 ;
    RECT -0.26 -0.27 0.26 0.27 ;
  LAYER bv3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER bm3 ;
    RECT -0.27 -0.27 0.27 0.27 ;
END BV3_400x400_540V_540H

VIA BV3_400x400_540V_540V
  LAYER bm4 ;
    RECT -0.27 -0.26 0.27 0.26 ;
  LAYER bv3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER bm3 ;
    RECT -0.27 -0.27 0.27 0.27 ;
END BV3_400x400_540V_540V

VIA BV3_400x400_540V_720d5H
  LAYER bm4 ;
    RECT -0.285 -0.36 0.285 0.36 ;
  LAYER bv3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER bm3 ;
    RECT -0.27 -0.27 0.27 0.27 ;
END BV3_400x400_540V_720d5H

VIA BV3_400x400_540V_720d5V
  LAYER bm4 ;
    RECT -0.36 -0.285 0.36 0.285 ;
  LAYER bv3 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER bm3 ;
    RECT -0.27 -0.27 0.27 0.27 ;
END BV3_400x400_540V_720d5V

VIA BV3_400x600_600V_1200d5H
  LAYER bm4 ;
    RECT -0.32 -0.6 0.32 0.6 ;
  LAYER bv3 ;
    RECT -0.2 -0.3 0.2 0.3 ;
  LAYER bm3 ;
    RECT -0.3 -0.4 0.3 0.4 ;
END BV3_400x600_600V_1200d5H

VIA BV3_400x600_600V_1200d5V
  LAYER bm4 ;
    RECT -0.6 -0.42 0.6 0.42 ;
  LAYER bv3 ;
    RECT -0.2 -0.3 0.2 0.3 ;
  LAYER bm3 ;
    RECT -0.3 -0.4 0.3 0.4 ;
END BV3_400x600_600V_1200d5V

VIA BV3_400x600_600V_2400d5H
  LAYER bm4 ;
    RECT -0.37 -1.2 0.37 1.2 ;
  LAYER bv3 ;
    RECT -0.2 -0.3 0.2 0.3 ;
  LAYER bm3 ;
    RECT -0.3 -0.4 0.3 0.4 ;
END BV3_400x600_600V_2400d5H

VIA BV3_400x600_600V_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.47 1.2 0.47 ;
  LAYER bv3 ;
    RECT -0.2 -0.3 0.2 0.3 ;
  LAYER bm3 ;
    RECT -0.3 -0.4 0.3 0.4 ;
END BV3_400x600_600V_2400d5V

VIA BV3_400x600_600V_540V
  LAYER bm4 ;
    RECT -0.27 -0.36 0.27 0.36 ;
  LAYER bv3 ;
    RECT -0.2 -0.3 0.2 0.3 ;
  LAYER bm3 ;
    RECT -0.3 -0.4 0.3 0.4 ;
END BV3_400x600_600V_540V

VIA BV3_400x600_600V_720H
  LAYER bm4 ;
    RECT -0.26 -0.36 0.26 0.36 ;
  LAYER bv3 ;
    RECT -0.2 -0.3 0.2 0.3 ;
  LAYER bm3 ;
    RECT -0.3 -0.4 0.3 0.4 ;
END BV3_400x600_600V_720H

VIA BV3_400x600_600V_720d5V
  LAYER bm4 ;
    RECT -0.36 -0.385 0.36 0.385 ;
  LAYER bv3 ;
    RECT -0.2 -0.3 0.2 0.3 ;
  LAYER bm3 ;
    RECT -0.3 -0.4 0.3 0.4 ;
END BV3_400x600_600V_720d5V

VIA BV3_400x600_600V_770H
  LAYER bm4 ;
    RECT -0.285 -0.385 0.285 0.385 ;
  LAYER bv3 ;
    RECT -0.2 -0.3 0.2 0.3 ;
  LAYER bm3 ;
    RECT -0.3 -0.4 0.3 0.4 ;
END BV3_400x600_600V_770H

VIA BV3_400x600_800H_1200d5H
  LAYER bm4 ;
    RECT -0.32 -0.6 0.32 0.6 ;
  LAYER bv3 ;
    RECT -0.2 -0.3 0.2 0.3 ;
  LAYER bm3 ;
    RECT -0.3 -0.4 0.3 0.4 ;
END BV3_400x600_800H_1200d5H

VIA BV3_400x600_800H_1200d5V
  LAYER bm4 ;
    RECT -0.6 -0.42 0.6 0.42 ;
  LAYER bv3 ;
    RECT -0.2 -0.3 0.2 0.3 ;
  LAYER bm3 ;
    RECT -0.3 -0.4 0.3 0.4 ;
END BV3_400x600_800H_1200d5V

VIA BV3_400x600_800H_2400d5H
  LAYER bm4 ;
    RECT -0.37 -1.2 0.37 1.2 ;
  LAYER bv3 ;
    RECT -0.2 -0.3 0.2 0.3 ;
  LAYER bm3 ;
    RECT -0.3 -0.4 0.3 0.4 ;
END BV3_400x600_800H_2400d5H

VIA BV3_400x600_800H_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.47 1.2 0.47 ;
  LAYER bv3 ;
    RECT -0.2 -0.3 0.2 0.3 ;
  LAYER bm3 ;
    RECT -0.3 -0.4 0.3 0.4 ;
END BV3_400x600_800H_2400d5V

VIA BV3_400x600_800H_540V
  LAYER bm4 ;
    RECT -0.27 -0.36 0.27 0.36 ;
  LAYER bv3 ;
    RECT -0.2 -0.3 0.2 0.3 ;
  LAYER bm3 ;
    RECT -0.3 -0.4 0.3 0.4 ;
END BV3_400x600_800H_540V

VIA BV3_400x600_800H_720H
  LAYER bm4 ;
    RECT -0.26 -0.36 0.26 0.36 ;
  LAYER bv3 ;
    RECT -0.2 -0.3 0.2 0.3 ;
  LAYER bm3 ;
    RECT -0.3 -0.4 0.3 0.4 ;
END BV3_400x600_800H_720H

VIA BV3_400x600_800H_720d5V
  LAYER bm4 ;
    RECT -0.36 -0.385 0.36 0.385 ;
  LAYER bv3 ;
    RECT -0.2 -0.3 0.2 0.3 ;
  LAYER bm3 ;
    RECT -0.3 -0.4 0.3 0.4 ;
END BV3_400x600_800H_720d5V

VIA BV3_400x600_800H_770H
  LAYER bm4 ;
    RECT -0.285 -0.385 0.285 0.385 ;
  LAYER bv3 ;
    RECT -0.2 -0.3 0.2 0.3 ;
  LAYER bm3 ;
    RECT -0.3 -0.4 0.3 0.4 ;
END BV3_400x600_800H_770H

VIA BV3_400x900_1100H_1070H
  LAYER bm4 ;
    RECT -0.285 -0.535 0.285 0.535 ;
  LAYER bv3 ;
    RECT -0.2 -0.45 0.2 0.45 ;
  LAYER bm3 ;
    RECT -0.3 -0.55 0.3 0.55 ;
END BV3_400x900_1100H_1070H

VIA BV3_400x900_1100H_1200d5H
  LAYER bm4 ;
    RECT -0.32 -0.6 0.32 0.6 ;
  LAYER bv3 ;
    RECT -0.2 -0.45 0.2 0.45 ;
  LAYER bm3 ;
    RECT -0.3 -0.55 0.3 0.55 ;
END BV3_400x900_1100H_1200d5H

VIA BV3_400x900_1100H_1200d5V
  LAYER bm4 ;
    RECT -0.6 -0.57 0.6 0.57 ;
  LAYER bv3 ;
    RECT -0.2 -0.45 0.2 0.45 ;
  LAYER bm3 ;
    RECT -0.3 -0.55 0.3 0.55 ;
END BV3_400x900_1100H_1200d5V

VIA BV3_400x900_1100H_2400d5H
  LAYER bm4 ;
    RECT -0.37 -1.2 0.37 1.2 ;
  LAYER bv3 ;
    RECT -0.2 -0.45 0.2 0.45 ;
  LAYER bm3 ;
    RECT -0.3 -0.55 0.3 0.55 ;
END BV3_400x900_1100H_2400d5H

VIA BV3_400x900_1100H_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.62 1.2 0.62 ;
  LAYER bv3 ;
    RECT -0.2 -0.45 0.2 0.45 ;
  LAYER bm3 ;
    RECT -0.3 -0.55 0.3 0.55 ;
END BV3_400x900_1100H_2400d5V

VIA BV3_400x900_1100H_540V
  LAYER bm4 ;
    RECT -0.27 -0.51 0.27 0.51 ;
  LAYER bv3 ;
    RECT -0.2 -0.45 0.2 0.45 ;
  LAYER bm3 ;
    RECT -0.3 -0.55 0.3 0.55 ;
END BV3_400x900_1100H_540V

VIA BV3_400x900_1100H_720d5V
  LAYER bm4 ;
    RECT -0.36 -0.535 0.36 0.535 ;
  LAYER bv3 ;
    RECT -0.2 -0.45 0.2 0.45 ;
  LAYER bm3 ;
    RECT -0.3 -0.55 0.3 0.55 ;
END BV3_400x900_1100H_720d5V

VIA BV3_400x900_600V_1070H
  LAYER bm4 ;
    RECT -0.285 -0.535 0.285 0.535 ;
  LAYER bv3 ;
    RECT -0.2 -0.45 0.2 0.45 ;
  LAYER bm3 ;
    RECT -0.3 -0.55 0.3 0.55 ;
END BV3_400x900_600V_1070H

VIA BV3_400x900_600V_1200d5H
  LAYER bm4 ;
    RECT -0.32 -0.6 0.32 0.6 ;
  LAYER bv3 ;
    RECT -0.2 -0.45 0.2 0.45 ;
  LAYER bm3 ;
    RECT -0.3 -0.55 0.3 0.55 ;
END BV3_400x900_600V_1200d5H

VIA BV3_400x900_600V_1200d5V
  LAYER bm4 ;
    RECT -0.6 -0.57 0.6 0.57 ;
  LAYER bv3 ;
    RECT -0.2 -0.45 0.2 0.45 ;
  LAYER bm3 ;
    RECT -0.3 -0.55 0.3 0.55 ;
END BV3_400x900_600V_1200d5V

VIA BV3_400x900_600V_2400d5H
  LAYER bm4 ;
    RECT -0.37 -1.2 0.37 1.2 ;
  LAYER bv3 ;
    RECT -0.2 -0.45 0.2 0.45 ;
  LAYER bm3 ;
    RECT -0.3 -0.55 0.3 0.55 ;
END BV3_400x900_600V_2400d5H

VIA BV3_400x900_600V_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.62 1.2 0.62 ;
  LAYER bv3 ;
    RECT -0.2 -0.45 0.2 0.45 ;
  LAYER bm3 ;
    RECT -0.3 -0.55 0.3 0.55 ;
END BV3_400x900_600V_2400d5V

VIA BV3_400x900_600V_540V
  LAYER bm4 ;
    RECT -0.27 -0.51 0.27 0.51 ;
  LAYER bv3 ;
    RECT -0.2 -0.45 0.2 0.45 ;
  LAYER bm3 ;
    RECT -0.3 -0.55 0.3 0.55 ;
END BV3_400x900_600V_540V

VIA BV3_400x900_600V_720d5V
  LAYER bm4 ;
    RECT -0.36 -0.535 0.36 0.535 ;
  LAYER bv3 ;
    RECT -0.2 -0.45 0.2 0.45 ;
  LAYER bm3 ;
    RECT -0.3 -0.55 0.3 0.55 ;
END BV3_400x900_600V_720d5V

VIA BV3_600x400_600H_1200d5H
  LAYER bm4 ;
    RECT -0.42 -0.6 0.42 0.6 ;
  LAYER bv3 ;
    RECT -0.3 -0.2 0.3 0.2 ;
  LAYER bm3 ;
    RECT -0.4 -0.3 0.4 0.3 ;
END BV3_600x400_600H_1200d5H

VIA BV3_600x400_600H_1200d5V
  LAYER bm4 ;
    RECT -0.6 -0.32 0.6 0.32 ;
  LAYER bv3 ;
    RECT -0.3 -0.2 0.3 0.2 ;
  LAYER bm3 ;
    RECT -0.4 -0.3 0.4 0.3 ;
END BV3_600x400_600H_1200d5V

VIA BV3_600x400_600H_2400d5H
  LAYER bm4 ;
    RECT -0.47 -1.2 0.47 1.2 ;
  LAYER bv3 ;
    RECT -0.3 -0.2 0.3 0.2 ;
  LAYER bm3 ;
    RECT -0.4 -0.3 0.4 0.3 ;
END BV3_600x400_600H_2400d5H

VIA BV3_600x400_600H_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.37 1.2 0.37 ;
  LAYER bv3 ;
    RECT -0.3 -0.2 0.3 0.2 ;
  LAYER bm3 ;
    RECT -0.4 -0.3 0.4 0.3 ;
END BV3_600x400_600H_2400d5V

VIA BV3_600x400_600H_540H
  LAYER bm4 ;
    RECT -0.36 -0.27 0.36 0.27 ;
  LAYER bv3 ;
    RECT -0.3 -0.2 0.3 0.2 ;
  LAYER bm3 ;
    RECT -0.4 -0.3 0.4 0.3 ;
END BV3_600x400_600H_540H

VIA BV3_600x400_600H_720V
  LAYER bm4 ;
    RECT -0.36 -0.26 0.36 0.26 ;
  LAYER bv3 ;
    RECT -0.3 -0.2 0.3 0.2 ;
  LAYER bm3 ;
    RECT -0.4 -0.3 0.4 0.3 ;
END BV3_600x400_600H_720V

VIA BV3_600x400_600H_720d5H
  LAYER bm4 ;
    RECT -0.385 -0.36 0.385 0.36 ;
  LAYER bv3 ;
    RECT -0.3 -0.2 0.3 0.2 ;
  LAYER bm3 ;
    RECT -0.4 -0.3 0.4 0.3 ;
END BV3_600x400_600H_720d5H

VIA BV3_600x400_600H_770V
  LAYER bm4 ;
    RECT -0.385 -0.285 0.385 0.285 ;
  LAYER bv3 ;
    RECT -0.3 -0.2 0.3 0.2 ;
  LAYER bm3 ;
    RECT -0.4 -0.3 0.4 0.3 ;
END BV3_600x400_600H_770V

VIA BV3_600x400_800V_1200d5H
  LAYER bm4 ;
    RECT -0.42 -0.6 0.42 0.6 ;
  LAYER bv3 ;
    RECT -0.3 -0.2 0.3 0.2 ;
  LAYER bm3 ;
    RECT -0.4 -0.3 0.4 0.3 ;
END BV3_600x400_800V_1200d5H

VIA BV3_600x400_800V_1200d5V
  LAYER bm4 ;
    RECT -0.6 -0.32 0.6 0.32 ;
  LAYER bv3 ;
    RECT -0.3 -0.2 0.3 0.2 ;
  LAYER bm3 ;
    RECT -0.4 -0.3 0.4 0.3 ;
END BV3_600x400_800V_1200d5V

VIA BV3_600x400_800V_2400d5H
  LAYER bm4 ;
    RECT -0.47 -1.2 0.47 1.2 ;
  LAYER bv3 ;
    RECT -0.3 -0.2 0.3 0.2 ;
  LAYER bm3 ;
    RECT -0.4 -0.3 0.4 0.3 ;
END BV3_600x400_800V_2400d5H

VIA BV3_600x400_800V_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.37 1.2 0.37 ;
  LAYER bv3 ;
    RECT -0.3 -0.2 0.3 0.2 ;
  LAYER bm3 ;
    RECT -0.4 -0.3 0.4 0.3 ;
END BV3_600x400_800V_2400d5V

VIA BV3_600x400_800V_540H
  LAYER bm4 ;
    RECT -0.36 -0.27 0.36 0.27 ;
  LAYER bv3 ;
    RECT -0.3 -0.2 0.3 0.2 ;
  LAYER bm3 ;
    RECT -0.4 -0.3 0.4 0.3 ;
END BV3_600x400_800V_540H

VIA BV3_600x400_800V_720V
  LAYER bm4 ;
    RECT -0.36 -0.26 0.36 0.26 ;
  LAYER bv3 ;
    RECT -0.3 -0.2 0.3 0.2 ;
  LAYER bm3 ;
    RECT -0.4 -0.3 0.4 0.3 ;
END BV3_600x400_800V_720V

VIA BV3_600x400_800V_720d5H
  LAYER bm4 ;
    RECT -0.385 -0.36 0.385 0.36 ;
  LAYER bv3 ;
    RECT -0.3 -0.2 0.3 0.2 ;
  LAYER bm3 ;
    RECT -0.4 -0.3 0.4 0.3 ;
END BV3_600x400_800V_720d5H

VIA BV3_600x400_800V_770V
  LAYER bm4 ;
    RECT -0.385 -0.285 0.385 0.285 ;
  LAYER bv3 ;
    RECT -0.3 -0.2 0.3 0.2 ;
  LAYER bm3 ;
    RECT -0.4 -0.3 0.4 0.3 ;
END BV3_600x400_800V_770V

VIA BV3_900x400_1100V_1070V
  LAYER bm4 ;
    RECT -0.535 -0.285 0.535 0.285 ;
  LAYER bv3 ;
    RECT -0.45 -0.2 0.45 0.2 ;
  LAYER bm3 ;
    RECT -0.55 -0.3 0.55 0.3 ;
END BV3_900x400_1100V_1070V

VIA BV3_900x400_1100V_1200d5H
  LAYER bm4 ;
    RECT -0.57 -0.6 0.57 0.6 ;
  LAYER bv3 ;
    RECT -0.45 -0.2 0.45 0.2 ;
  LAYER bm3 ;
    RECT -0.55 -0.3 0.55 0.3 ;
END BV3_900x400_1100V_1200d5H

VIA BV3_900x400_1100V_1200d5V
  LAYER bm4 ;
    RECT -0.6 -0.32 0.6 0.32 ;
  LAYER bv3 ;
    RECT -0.45 -0.2 0.45 0.2 ;
  LAYER bm3 ;
    RECT -0.55 -0.3 0.55 0.3 ;
END BV3_900x400_1100V_1200d5V

VIA BV3_900x400_1100V_2400d5H
  LAYER bm4 ;
    RECT -0.62 -1.2 0.62 1.2 ;
  LAYER bv3 ;
    RECT -0.45 -0.2 0.45 0.2 ;
  LAYER bm3 ;
    RECT -0.55 -0.3 0.55 0.3 ;
END BV3_900x400_1100V_2400d5H

VIA BV3_900x400_1100V_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.37 1.2 0.37 ;
  LAYER bv3 ;
    RECT -0.45 -0.2 0.45 0.2 ;
  LAYER bm3 ;
    RECT -0.55 -0.3 0.55 0.3 ;
END BV3_900x400_1100V_2400d5V

VIA BV3_900x400_1100V_540H
  LAYER bm4 ;
    RECT -0.51 -0.27 0.51 0.27 ;
  LAYER bv3 ;
    RECT -0.45 -0.2 0.45 0.2 ;
  LAYER bm3 ;
    RECT -0.55 -0.3 0.55 0.3 ;
END BV3_900x400_1100V_540H

VIA BV3_900x400_1100V_720d5H
  LAYER bm4 ;
    RECT -0.535 -0.36 0.535 0.36 ;
  LAYER bv3 ;
    RECT -0.45 -0.2 0.45 0.2 ;
  LAYER bm3 ;
    RECT -0.55 -0.3 0.55 0.3 ;
END BV3_900x400_1100V_720d5H

VIA BV3_900x400_600H_1070V
  LAYER bm4 ;
    RECT -0.535 -0.285 0.535 0.285 ;
  LAYER bv3 ;
    RECT -0.45 -0.2 0.45 0.2 ;
  LAYER bm3 ;
    RECT -0.55 -0.3 0.55 0.3 ;
END BV3_900x400_600H_1070V

VIA BV3_900x400_600H_1200d5H
  LAYER bm4 ;
    RECT -0.57 -0.6 0.57 0.6 ;
  LAYER bv3 ;
    RECT -0.45 -0.2 0.45 0.2 ;
  LAYER bm3 ;
    RECT -0.55 -0.3 0.55 0.3 ;
END BV3_900x400_600H_1200d5H

VIA BV3_900x400_600H_1200d5V
  LAYER bm4 ;
    RECT -0.6 -0.32 0.6 0.32 ;
  LAYER bv3 ;
    RECT -0.45 -0.2 0.45 0.2 ;
  LAYER bm3 ;
    RECT -0.55 -0.3 0.55 0.3 ;
END BV3_900x400_600H_1200d5V

VIA BV3_900x400_600H_2400d5H
  LAYER bm4 ;
    RECT -0.62 -1.2 0.62 1.2 ;
  LAYER bv3 ;
    RECT -0.45 -0.2 0.45 0.2 ;
  LAYER bm3 ;
    RECT -0.55 -0.3 0.55 0.3 ;
END BV3_900x400_600H_2400d5H

VIA BV3_900x400_600H_2400d5V
  LAYER bm4 ;
    RECT -1.2 -0.37 1.2 0.37 ;
  LAYER bv3 ;
    RECT -0.45 -0.2 0.45 0.2 ;
  LAYER bm3 ;
    RECT -0.55 -0.3 0.55 0.3 ;
END BV3_900x400_600H_2400d5V

VIA BV3_900x400_600H_540H
  LAYER bm4 ;
    RECT -0.51 -0.27 0.51 0.27 ;
  LAYER bv3 ;
    RECT -0.45 -0.2 0.45 0.2 ;
  LAYER bm3 ;
    RECT -0.55 -0.3 0.55 0.3 ;
END BV3_900x400_600H_540H

VIA BV3_900x400_600H_720d5H
  LAYER bm4 ;
    RECT -0.535 -0.36 0.535 0.36 ;
  LAYER bv3 ;
    RECT -0.45 -0.2 0.45 0.2 ;
  LAYER bm3 ;
    RECT -0.55 -0.3 0.55 0.3 ;
END BV3_900x400_600H_720d5H

VIA BV4_1800x800_1080H_2000H
  LAYER bm5 ;
    RECT -1.5 -1 1.5 1 ;
  LAYER bv4 ;
    RECT -0.9 -0.4 0.9 0.4 ;
  LAYER bm4 ;
    RECT -1.04 -0.54 1.04 0.54 ;
END BV4_1800x800_1080H_2000H

VIA BV4_1800x800_1080H_3000V
  LAYER bm5 ;
    RECT -1.5 -1 1.5 1 ;
  LAYER bv4 ;
    RECT -0.9 -0.4 0.9 0.4 ;
  LAYER bm4 ;
    RECT -1.04 -0.54 1.04 0.54 ;
END BV4_1800x800_1080H_3000V

VIA BV4_1800x800_2080V_2000H
  LAYER bm5 ;
    RECT -1.5 -1 1.5 1 ;
  LAYER bv4 ;
    RECT -0.9 -0.4 0.9 0.4 ;
  LAYER bm4 ;
    RECT -1.04 -0.54 1.04 0.54 ;
END BV4_1800x800_2080V_2000H

VIA BV4_1800x800_2080V_3000V
  LAYER bm5 ;
    RECT -1.5 -1 1.5 1 ;
  LAYER bv4 ;
    RECT -0.9 -0.4 0.9 0.4 ;
  LAYER bm4 ;
    RECT -1.04 -0.54 1.04 0.54 ;
END BV4_1800x800_2080V_3000V

VIA BV4_1850x800_1080H_2000H
  LAYER bm5 ;
    RECT -1.525 -1 1.525 1 ;
  LAYER bv4 ;
    RECT -0.925 -0.4 0.925 0.4 ;
  LAYER bm4 ;
    RECT -1.065 -0.54 1.065 0.54 ;
END BV4_1850x800_1080H_2000H

VIA BV4_1850x800_1080H_3050V
  LAYER bm5 ;
    RECT -1.525 -1 1.525 1 ;
  LAYER bv4 ;
    RECT -0.925 -0.4 0.925 0.4 ;
  LAYER bm4 ;
    RECT -1.065 -0.54 1.065 0.54 ;
END BV4_1850x800_1080H_3050V

VIA BV4_1850x800_2130V_2000H
  LAYER bm5 ;
    RECT -1.525 -1 1.525 1 ;
  LAYER bv4 ;
    RECT -0.925 -0.4 0.925 0.4 ;
  LAYER bm4 ;
    RECT -1.065 -0.54 1.065 0.54 ;
END BV4_1850x800_2130V_2000H

VIA BV4_1850x800_2130V_3050V
  LAYER bm5 ;
    RECT -1.525 -1 1.525 1 ;
  LAYER bv4 ;
    RECT -0.925 -0.4 0.925 0.4 ;
  LAYER bm4 ;
    RECT -1.065 -0.54 1.065 0.54 ;
END BV4_1850x800_2130V_3050V

VIA BV4_2800x800_1080H_2000H
  LAYER bm5 ;
    RECT -2 -1 2 1 ;
  LAYER bv4 ;
    RECT -1.4 -0.4 1.4 0.4 ;
  LAYER bm4 ;
    RECT -1.54 -0.54 1.54 0.54 ;
END BV4_2800x800_1080H_2000H

VIA BV4_2800x800_1080H_4000V
  LAYER bm5 ;
    RECT -2 -1 2 1 ;
  LAYER bv4 ;
    RECT -1.4 -0.4 1.4 0.4 ;
  LAYER bm4 ;
    RECT -1.54 -0.54 1.54 0.54 ;
END BV4_2800x800_1080H_4000V

VIA BV4_2800x800_3080V_2000H
  LAYER bm5 ;
    RECT -2 -1 2 1 ;
  LAYER bv4 ;
    RECT -1.4 -0.4 1.4 0.4 ;
  LAYER bm4 ;
    RECT -1.54 -0.54 1.54 0.54 ;
END BV4_2800x800_3080V_2000H

VIA BV4_2800x800_3080V_4000V
  LAYER bm5 ;
    RECT -2 -1 2 1 ;
  LAYER bv4 ;
    RECT -1.4 -0.4 1.4 0.4 ;
  LAYER bm4 ;
    RECT -1.54 -0.54 1.54 0.54 ;
END BV4_2800x800_3080V_4000V

VIA BV4_3700x800_1080H_2000H
  LAYER bm5 ;
    RECT -2.45 -1 2.45 1 ;
  LAYER bv4 ;
    RECT -1.85 -0.4 1.85 0.4 ;
  LAYER bm4 ;
    RECT -1.99 -0.54 1.99 0.54 ;
END BV4_3700x800_1080H_2000H

VIA BV4_3700x800_1080H_4900V
  LAYER bm5 ;
    RECT -2.45 -1 2.45 1 ;
  LAYER bv4 ;
    RECT -1.85 -0.4 1.85 0.4 ;
  LAYER bm4 ;
    RECT -1.99 -0.54 1.99 0.54 ;
END BV4_3700x800_1080H_4900V

VIA BV4_3700x800_3980V_2000H
  LAYER bm5 ;
    RECT -2.45 -1 2.45 1 ;
  LAYER bv4 ;
    RECT -1.85 -0.4 1.85 0.4 ;
  LAYER bm4 ;
    RECT -1.99 -0.54 1.99 0.54 ;
END BV4_3700x800_3980V_2000H

VIA BV4_3700x800_3980V_4900V
  LAYER bm5 ;
    RECT -2.45 -1 2.45 1 ;
  LAYER bv4 ;
    RECT -1.85 -0.4 1.85 0.4 ;
  LAYER bm4 ;
    RECT -1.99 -0.54 1.99 0.54 ;
END BV4_3700x800_3980V_4900V

VIA BV4_5000x800_1080H_2000H
  LAYER bm5 ;
    RECT -3.1 -1 3.1 1 ;
  LAYER bv4 ;
    RECT -2.5 -0.4 2.5 0.4 ;
  LAYER bm4 ;
    RECT -2.64 -0.54 2.64 0.54 ;
END BV4_5000x800_1080H_2000H

VIA BV4_5000x800_1080H_6200V
  LAYER bm5 ;
    RECT -3.1 -1 3.1 1 ;
  LAYER bv4 ;
    RECT -2.5 -0.4 2.5 0.4 ;
  LAYER bm4 ;
    RECT -2.64 -0.54 2.64 0.54 ;
END BV4_5000x800_1080H_6200V

VIA BV4_5000x800_5280V_2000H
  LAYER bm5 ;
    RECT -3.1 -1 3.1 1 ;
  LAYER bv4 ;
    RECT -2.5 -0.4 2.5 0.4 ;
  LAYER bm4 ;
    RECT -2.64 -0.54 2.64 0.54 ;
END BV4_5000x800_5280V_2000H

VIA BV4_5000x800_5280V_6200V
  LAYER bm5 ;
    RECT -3.1 -1 3.1 1 ;
  LAYER bv4 ;
    RECT -2.5 -0.4 2.5 0.4 ;
  LAYER bm4 ;
    RECT -2.64 -0.54 2.64 0.54 ;
END BV4_5000x800_5280V_6200V

VIA BV4_7400x800_1080H_2000H
  LAYER bm5 ;
    RECT -4.3 -1 4.3 1 ;
  LAYER bv4 ;
    RECT -3.7 -0.4 3.7 0.4 ;
  LAYER bm4 ;
    RECT -3.84 -0.54 3.84 0.54 ;
END BV4_7400x800_1080H_2000H

VIA BV4_7400x800_1080H_8600V
  LAYER bm5 ;
    RECT -4.3 -1 4.3 1 ;
  LAYER bv4 ;
    RECT -3.7 -0.4 3.7 0.4 ;
  LAYER bm4 ;
    RECT -3.84 -0.54 3.84 0.54 ;
END BV4_7400x800_1080H_8600V

VIA BV4_800x1800_1080V_2000V
  LAYER bm5 ;
    RECT -1 -1.5 1 1.5 ;
  LAYER bv4 ;
    RECT -0.4 -0.9 0.4 0.9 ;
  LAYER bm4 ;
    RECT -0.54 -1.04 0.54 1.04 ;
END BV4_800x1800_1080V_2000V

VIA BV4_800x1800_1080V_3000H
  LAYER bm5 ;
    RECT -1 -1.5 1 1.5 ;
  LAYER bv4 ;
    RECT -0.4 -0.9 0.4 0.9 ;
  LAYER bm4 ;
    RECT -0.54 -1.04 0.54 1.04 ;
END BV4_800x1800_1080V_3000H

VIA BV4_800x1800_2080H_2000V
  LAYER bm5 ;
    RECT -1 -1.5 1 1.5 ;
  LAYER bv4 ;
    RECT -0.4 -0.9 0.4 0.9 ;
  LAYER bm4 ;
    RECT -0.54 -1.04 0.54 1.04 ;
END BV4_800x1800_2080H_2000V

VIA BV4_800x1800_2080H_3000H
  LAYER bm5 ;
    RECT -1 -1.5 1 1.5 ;
  LAYER bv4 ;
    RECT -0.4 -0.9 0.4 0.9 ;
  LAYER bm4 ;
    RECT -0.54 -1.04 0.54 1.04 ;
END BV4_800x1800_2080H_3000H

VIA BV4_800x1850_1080V_2000V
  LAYER bm5 ;
    RECT -1 -1.525 1 1.525 ;
  LAYER bv4 ;
    RECT -0.4 -0.925 0.4 0.925 ;
  LAYER bm4 ;
    RECT -0.54 -1.065 0.54 1.065 ;
END BV4_800x1850_1080V_2000V

VIA BV4_800x1850_1080V_3050H
  LAYER bm5 ;
    RECT -1 -1.525 1 1.525 ;
  LAYER bv4 ;
    RECT -0.4 -0.925 0.4 0.925 ;
  LAYER bm4 ;
    RECT -0.54 -1.065 0.54 1.065 ;
END BV4_800x1850_1080V_3050H

VIA BV4_800x1850_2130H_2000V
  LAYER bm5 ;
    RECT -1 -1.525 1 1.525 ;
  LAYER bv4 ;
    RECT -0.4 -0.925 0.4 0.925 ;
  LAYER bm4 ;
    RECT -0.54 -1.065 0.54 1.065 ;
END BV4_800x1850_2130H_2000V

VIA BV4_800x1850_2130H_3050H
  LAYER bm5 ;
    RECT -1 -1.525 1 1.525 ;
  LAYER bv4 ;
    RECT -0.4 -0.925 0.4 0.925 ;
  LAYER bm4 ;
    RECT -0.54 -1.065 0.54 1.065 ;
END BV4_800x1850_2130H_3050H

VIA BV4_800x2800_1080V_2000V
  LAYER bm5 ;
    RECT -1 -2 1 2 ;
  LAYER bv4 ;
    RECT -0.4 -1.4 0.4 1.4 ;
  LAYER bm4 ;
    RECT -0.54 -1.54 0.54 1.54 ;
END BV4_800x2800_1080V_2000V

VIA BV4_800x2800_1080V_4000H
  LAYER bm5 ;
    RECT -1 -2 1 2 ;
  LAYER bv4 ;
    RECT -0.4 -1.4 0.4 1.4 ;
  LAYER bm4 ;
    RECT -0.54 -1.54 0.54 1.54 ;
END BV4_800x2800_1080V_4000H

VIA BV4_800x2800_3080H_2000V
  LAYER bm5 ;
    RECT -1 -2 1 2 ;
  LAYER bv4 ;
    RECT -0.4 -1.4 0.4 1.4 ;
  LAYER bm4 ;
    RECT -0.54 -1.54 0.54 1.54 ;
END BV4_800x2800_3080H_2000V

VIA BV4_800x2800_3080H_4000H
  LAYER bm5 ;
    RECT -1 -2 1 2 ;
  LAYER bv4 ;
    RECT -0.4 -1.4 0.4 1.4 ;
  LAYER bm4 ;
    RECT -0.54 -1.54 0.54 1.54 ;
END BV4_800x2800_3080H_4000H

VIA BV4_800x3700_1080V_2000V
  LAYER bm5 ;
    RECT -1 -2.45 1 2.45 ;
  LAYER bv4 ;
    RECT -0.4 -1.85 0.4 1.85 ;
  LAYER bm4 ;
    RECT -0.54 -1.99 0.54 1.99 ;
END BV4_800x3700_1080V_2000V

VIA BV4_800x3700_1080V_4900H
  LAYER bm5 ;
    RECT -1 -2.45 1 2.45 ;
  LAYER bv4 ;
    RECT -0.4 -1.85 0.4 1.85 ;
  LAYER bm4 ;
    RECT -0.54 -1.99 0.54 1.99 ;
END BV4_800x3700_1080V_4900H

VIA BV4_800x3700_3980H_2000V
  LAYER bm5 ;
    RECT -1 -2.45 1 2.45 ;
  LAYER bv4 ;
    RECT -0.4 -1.85 0.4 1.85 ;
  LAYER bm4 ;
    RECT -0.54 -1.99 0.54 1.99 ;
END BV4_800x3700_3980H_2000V

VIA BV4_800x3700_3980H_4900H
  LAYER bm5 ;
    RECT -1 -2.45 1 2.45 ;
  LAYER bv4 ;
    RECT -0.4 -1.85 0.4 1.85 ;
  LAYER bm4 ;
    RECT -0.54 -1.99 0.54 1.99 ;
END BV4_800x3700_3980H_4900H

VIA BV4_800x5000_1080V_2000V
  LAYER bm5 ;
    RECT -1 -3.1 1 3.1 ;
  LAYER bv4 ;
    RECT -0.4 -2.5 0.4 2.5 ;
  LAYER bm4 ;
    RECT -0.54 -2.64 0.54 2.64 ;
END BV4_800x5000_1080V_2000V

VIA BV4_800x5000_1080V_6200H
  LAYER bm5 ;
    RECT -1 -3.1 1 3.1 ;
  LAYER bv4 ;
    RECT -0.4 -2.5 0.4 2.5 ;
  LAYER bm4 ;
    RECT -0.54 -2.64 0.54 2.64 ;
END BV4_800x5000_1080V_6200H

VIA BV4_800x5000_5280H_2000V
  LAYER bm5 ;
    RECT -1 -3.1 1 3.1 ;
  LAYER bv4 ;
    RECT -0.4 -2.5 0.4 2.5 ;
  LAYER bm4 ;
    RECT -0.54 -2.64 0.54 2.64 ;
END BV4_800x5000_5280H_2000V

VIA BV4_800x5000_5280H_6200H
  LAYER bm5 ;
    RECT -1 -3.1 1 3.1 ;
  LAYER bv4 ;
    RECT -0.4 -2.5 0.4 2.5 ;
  LAYER bm4 ;
    RECT -0.54 -2.64 0.54 2.64 ;
END BV4_800x5000_5280H_6200H

VIA BV4_800x7400_1080V_2000V
  LAYER bm5 ;
    RECT -1 -4.3 1 4.3 ;
  LAYER bv4 ;
    RECT -0.4 -3.7 0.4 3.7 ;
  LAYER bm4 ;
    RECT -0.54 -3.84 0.54 3.84 ;
END BV4_800x7400_1080V_2000V

VIA BV4_800x7400_1080V_8600H
  LAYER bm5 ;
    RECT -1 -4.3 1 4.3 ;
  LAYER bv4 ;
    RECT -0.4 -3.7 0.4 3.7 ;
  LAYER bm4 ;
    RECT -0.54 -3.84 0.54 3.84 ;
END BV4_800x7400_1080V_8600H

VIA V0_30x20_20H_30V
  LAYER m0 ;
    RECT -0.017 -0.01 0.017 0.01 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.015 -0.021 0.015 0.021 ;
END V0_30x20_20H_30V

VIA V0_30x20_20H_35H
  LAYER m0 ;
    RECT -0.017 -0.01 0.017 0.01 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.026 -0.0175 0.026 0.0175 ;
END V0_30x20_20H_35H

VIA V0_30x20_20H_56H
  LAYER m0 ;
    RECT -0.017 -0.01 0.017 0.01 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.026 -0.028 0.026 0.028 ;
END V0_30x20_20H_56H

VIA V0_30x20_20H_56V
  LAYER m0 ;
    RECT -0.017 -0.01 0.017 0.01 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.028 -0.021 0.028 0.021 ;
END V0_30x20_20H_56V

VIA V0_30x20_20H_70V
  LAYER m0 ;
    RECT -0.017 -0.01 0.017 0.01 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.035 -0.021 0.035 0.021 ;
END V0_30x20_20H_70V

VIA V0_30x20_28H_30V
  LAYER m0 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.015 -0.021 0.015 0.021 ;
END V0_30x20_28H_30V

VIA V0_30x20_28H_35H
  LAYER m0 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.026 -0.0175 0.026 0.0175 ;
END V0_30x20_28H_35H

VIA V0_30x20_28H_56H
  LAYER m0 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.026 -0.028 0.026 0.028 ;
END V0_30x20_28H_56H

VIA V0_30x20_28H_56V
  LAYER m0 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.028 -0.021 0.028 0.021 ;
END V0_30x20_28H_56V

VIA V0_30x20_28H_70V
  LAYER m0 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.035 -0.021 0.035 0.021 ;
END V0_30x20_28H_70V

VIA V0_30x20_38H_30V
  LAYER m0 ;
    RECT -0.017 -0.019 0.017 0.019 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.015 -0.021 0.015 0.021 ;
END V0_30x20_38H_30V

VIA V0_30x20_38H_35H
  LAYER m0 ;
    RECT -0.017 -0.019 0.017 0.019 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.026 -0.0175 0.026 0.0175 ;
END V0_30x20_38H_35H

VIA V0_30x20_38H_56H
  LAYER m0 ;
    RECT -0.017 -0.019 0.017 0.019 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.026 -0.028 0.026 0.028 ;
END V0_30x20_38H_56H

VIA V0_30x20_38H_56V
  LAYER m0 ;
    RECT -0.017 -0.019 0.017 0.019 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.028 -0.021 0.028 0.021 ;
END V0_30x20_38H_56V

VIA V0_30x20_38H_70V
  LAYER m0 ;
    RECT -0.017 -0.019 0.017 0.019 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.035 -0.021 0.035 0.021 ;
END V0_30x20_38H_70V

VIA V0_30x20_56H_30V
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.015 -0.021 0.015 0.021 ;
END V0_30x20_56H_30V

VIA V0_30x20_56H_35H
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.026 -0.0175 0.026 0.0175 ;
END V0_30x20_56H_35H

VIA V0_30x20_56H_56H
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.026 -0.028 0.026 0.028 ;
END V0_30x20_56H_56H

VIA V0_30x20_56H_56V
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.028 -0.021 0.028 0.021 ;
END V0_30x20_56H_56V

VIA V0_30x20_56H_70V
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m1 ;
    RECT -0.035 -0.021 0.035 0.021 ;
END V0_30x20_56H_70V

VIA V0_30x28_28H_30V
  LAYER m0 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER v0 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m1 ;
    RECT -0.015 -0.025 0.015 0.025 ;
END V0_30x28_28H_30V

VIA V0_30x28_28H_35H
  LAYER m0 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER v0 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m1 ;
    RECT -0.026 -0.0175 0.026 0.0175 ;
END V0_30x28_28H_35H

VIA V0_30x28_28H_56H
  LAYER m0 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER v0 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m1 ;
    RECT -0.026 -0.028 0.026 0.028 ;
END V0_30x28_28H_56H

VIA V0_30x28_28H_56V
  LAYER m0 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER v0 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m1 ;
    RECT -0.028 -0.025 0.028 0.025 ;
END V0_30x28_28H_56V

VIA V0_30x28_28H_70V
  LAYER m0 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER v0 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m1 ;
    RECT -0.035 -0.025 0.035 0.025 ;
END V0_30x28_28H_70V

VIA V0_30x28_38H_30V
  LAYER m0 ;
    RECT -0.017 -0.019 0.017 0.019 ;
  LAYER v0 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m1 ;
    RECT -0.015 -0.025 0.015 0.025 ;
END V0_30x28_38H_30V

VIA V0_30x28_38H_35H
  LAYER m0 ;
    RECT -0.017 -0.019 0.017 0.019 ;
  LAYER v0 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m1 ;
    RECT -0.026 -0.0175 0.026 0.0175 ;
END V0_30x28_38H_35H

VIA V0_30x28_38H_56H
  LAYER m0 ;
    RECT -0.017 -0.019 0.017 0.019 ;
  LAYER v0 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m1 ;
    RECT -0.026 -0.028 0.026 0.028 ;
END V0_30x28_38H_56H

VIA V0_30x28_38H_56V
  LAYER m0 ;
    RECT -0.017 -0.019 0.017 0.019 ;
  LAYER v0 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m1 ;
    RECT -0.028 -0.025 0.028 0.025 ;
END V0_30x28_38H_56V

VIA V0_30x28_38H_70V
  LAYER m0 ;
    RECT -0.017 -0.019 0.017 0.019 ;
  LAYER v0 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m1 ;
    RECT -0.035 -0.025 0.035 0.025 ;
END V0_30x28_38H_70V

VIA V0_30x28_56H_30V
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m1 ;
    RECT -0.015 -0.025 0.015 0.025 ;
END V0_30x28_56H_30V

VIA V0_30x28_56H_35H
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m1 ;
    RECT -0.026 -0.0175 0.026 0.0175 ;
END V0_30x28_56H_35H

VIA V0_30x28_56H_56H
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m1 ;
    RECT -0.026 -0.028 0.026 0.028 ;
END V0_30x28_56H_56H

VIA V0_30x28_56H_56V
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m1 ;
    RECT -0.028 -0.025 0.028 0.025 ;
END V0_30x28_56H_56V

VIA V0_30x28_56H_70V
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m1 ;
    RECT -0.035 -0.025 0.035 0.025 ;
END V0_30x28_56H_70V

VIA V0_30x38_38H_30V
  LAYER m0 ;
    RECT -0.017 -0.019 0.017 0.019 ;
  LAYER v0 ;
    RECT -0.015 -0.019 0.015 0.019 ;
  LAYER m1 ;
    RECT -0.015 -0.03 0.015 0.03 ;
END V0_30x38_38H_30V

VIA V0_30x38_38H_56H
  LAYER m0 ;
    RECT -0.017 -0.019 0.017 0.019 ;
  LAYER v0 ;
    RECT -0.015 -0.019 0.015 0.019 ;
  LAYER m1 ;
    RECT -0.026 -0.028 0.026 0.028 ;
END V0_30x38_38H_56H

VIA V0_30x38_38H_56V
  LAYER m0 ;
    RECT -0.017 -0.019 0.017 0.019 ;
  LAYER v0 ;
    RECT -0.015 -0.019 0.015 0.019 ;
  LAYER m1 ;
    RECT -0.028 -0.03 0.028 0.03 ;
END V0_30x38_38H_56V

VIA V0_30x38_38H_70V
  LAYER m0 ;
    RECT -0.017 -0.019 0.017 0.019 ;
  LAYER v0 ;
    RECT -0.015 -0.019 0.015 0.019 ;
  LAYER m1 ;
    RECT -0.035 -0.03 0.035 0.03 ;
END V0_30x38_38H_70V

VIA V0_30x38_56H_30V
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.019 0.015 0.019 ;
  LAYER m1 ;
    RECT -0.015 -0.03 0.015 0.03 ;
END V0_30x38_56H_30V

VIA V0_30x38_56H_56H
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.019 0.015 0.019 ;
  LAYER m1 ;
    RECT -0.026 -0.028 0.026 0.028 ;
END V0_30x38_56H_56H

VIA V0_30x38_56H_56V
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.019 0.015 0.019 ;
  LAYER m1 ;
    RECT -0.028 -0.03 0.028 0.03 ;
END V0_30x38_56H_56V

VIA V0_30x38_56H_70V
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.019 0.015 0.019 ;
  LAYER m1 ;
    RECT -0.035 -0.03 0.035 0.03 ;
END V0_30x38_56H_70V

VIA V0_30x56B_20H_30V
  LAYER m0 ;
    RECT -0.017 -0.01 0.017 0.01 ;
  LAYER v0 ;
    RECT -0.015 -0.028 0.015 0.028 ;
  LAYER m1 ;
    RECT -0.015 -0.033 0.015 0.033 ;
END V0_30x56B_20H_30V

VIA V0_30x56B_20H_56H
  LAYER m0 ;
    RECT -0.017 -0.01 0.017 0.01 ;
  LAYER v0 ;
    RECT -0.015 -0.028 0.015 0.028 ;
  LAYER m1 ;
    RECT -0.026 -0.028 0.026 0.028 ;
END V0_30x56B_20H_56H

VIA V0_30x56B_20H_56V
  LAYER m0 ;
    RECT -0.017 -0.01 0.017 0.01 ;
  LAYER v0 ;
    RECT -0.015 -0.028 0.015 0.028 ;
  LAYER m1 ;
    RECT -0.028 -0.033 0.028 0.033 ;
END V0_30x56B_20H_56V

VIA V0_30x56B_20H_70V
  LAYER m0 ;
    RECT -0.017 -0.01 0.017 0.01 ;
  LAYER v0 ;
    RECT -0.015 -0.028 0.015 0.028 ;
  LAYER m1 ;
    RECT -0.035 -0.033 0.035 0.033 ;
END V0_30x56B_20H_70V

VIA V0_30x56_56H_30V
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.028 0.015 0.028 ;
  LAYER m1 ;
    RECT -0.015 -0.033 0.015 0.033 ;
END V0_30x56_56H_30V

VIA V0_30x56_56H_56H
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.028 0.015 0.028 ;
  LAYER m1 ;
    RECT -0.026 -0.028 0.026 0.028 ;
END V0_30x56_56H_56H

VIA V0_30x56_56H_56V
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.028 0.015 0.028 ;
  LAYER m1 ;
    RECT -0.028 -0.033 0.028 0.033 ;
END V0_30x56_56H_56V

VIA V0_30x56_56H_70V
  LAYER m0 ;
    RECT -0.017 -0.028 0.017 0.028 ;
  LAYER v0 ;
    RECT -0.015 -0.028 0.015 0.028 ;
  LAYER m1 ;
    RECT -0.035 -0.033 0.035 0.033 ;
END V0_30x56_56H_70V

VIA V0_35x35_38H_35H
  LAYER m0 ;
    RECT -0.0195 -0.019 0.0195 0.019 ;
  LAYER v0 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m1 ;
    RECT -0.0225 -0.0175 0.0225 0.0175 ;
END V0_35x35_38H_35H

VIA V0_35x35_38H_56H
  LAYER m0 ;
    RECT -0.0195 -0.019 0.0195 0.019 ;
  LAYER v0 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m1 ;
    RECT -0.0225 -0.028 0.0225 0.028 ;
END V0_35x35_38H_56H

VIA V0_35x35_38H_56V
  LAYER m0 ;
    RECT -0.0195 -0.019 0.0195 0.019 ;
  LAYER v0 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m1 ;
    RECT -0.028 -0.0225 0.028 0.0225 ;
END V0_35x35_38H_56V

VIA V0_35x35_38H_70V
  LAYER m0 ;
    RECT -0.0195 -0.019 0.0195 0.019 ;
  LAYER v0 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m1 ;
    RECT -0.035 -0.0225 0.035 0.0225 ;
END V0_35x35_38H_70V

VIA V0_35x35_56H_35H
  LAYER m0 ;
    RECT -0.0195 -0.028 0.0195 0.028 ;
  LAYER v0 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m1 ;
    RECT -0.0225 -0.0175 0.0225 0.0175 ;
END V0_35x35_56H_35H

VIA V0_35x35_56H_56H
  LAYER m0 ;
    RECT -0.0195 -0.028 0.0195 0.028 ;
  LAYER v0 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m1 ;
    RECT -0.0225 -0.028 0.0225 0.028 ;
END V0_35x35_56H_56H

VIA V0_35x35_56H_56V
  LAYER m0 ;
    RECT -0.0195 -0.028 0.0195 0.028 ;
  LAYER v0 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m1 ;
    RECT -0.028 -0.0225 0.028 0.0225 ;
END V0_35x35_56H_56V

VIA V0_35x35_56H_70V
  LAYER m0 ;
    RECT -0.0195 -0.028 0.0195 0.028 ;
  LAYER v0 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m1 ;
    RECT -0.035 -0.0225 0.035 0.0225 ;
END V0_35x35_56H_70V

VIA V0_56x20_20H_35H
  LAYER m0 ;
    RECT -0.03 -0.01 0.03 0.01 ;
  LAYER v0 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m1 ;
    RECT -0.039 -0.0175 0.039 0.0175 ;
END V0_56x20_20H_35H

VIA V0_56x20_20H_56H
  LAYER m0 ;
    RECT -0.03 -0.01 0.03 0.01 ;
  LAYER v0 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m1 ;
    RECT -0.039 -0.028 0.039 0.028 ;
END V0_56x20_20H_56H

VIA V0_56x20_20H_56V
  LAYER m0 ;
    RECT -0.03 -0.01 0.03 0.01 ;
  LAYER v0 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m1 ;
    RECT -0.028 -0.021 0.028 0.021 ;
END V0_56x20_20H_56V

VIA V0_56x20_20H_70V
  LAYER m0 ;
    RECT -0.03 -0.01 0.03 0.01 ;
  LAYER v0 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m1 ;
    RECT -0.035 -0.021 0.035 0.021 ;
END V0_56x20_20H_70V

VIA V0_56x20_28H_35H
  LAYER m0 ;
    RECT -0.03 -0.014 0.03 0.014 ;
  LAYER v0 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m1 ;
    RECT -0.039 -0.0175 0.039 0.0175 ;
END V0_56x20_28H_35H

VIA V0_56x20_28H_56H
  LAYER m0 ;
    RECT -0.03 -0.014 0.03 0.014 ;
  LAYER v0 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m1 ;
    RECT -0.039 -0.028 0.039 0.028 ;
END V0_56x20_28H_56H

VIA V0_56x20_28H_56V
  LAYER m0 ;
    RECT -0.03 -0.014 0.03 0.014 ;
  LAYER v0 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m1 ;
    RECT -0.028 -0.021 0.028 0.021 ;
END V0_56x20_28H_56V

VIA V0_56x20_28H_70V
  LAYER m0 ;
    RECT -0.03 -0.014 0.03 0.014 ;
  LAYER v0 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m1 ;
    RECT -0.035 -0.021 0.035 0.021 ;
END V0_56x20_28H_70V

VIA V0_56x20_38H_35H
  LAYER m0 ;
    RECT -0.03 -0.019 0.03 0.019 ;
  LAYER v0 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m1 ;
    RECT -0.039 -0.0175 0.039 0.0175 ;
END V0_56x20_38H_35H

VIA V0_56x20_38H_56H
  LAYER m0 ;
    RECT -0.03 -0.019 0.03 0.019 ;
  LAYER v0 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m1 ;
    RECT -0.039 -0.028 0.039 0.028 ;
END V0_56x20_38H_56H

VIA V0_56x20_38H_56V
  LAYER m0 ;
    RECT -0.03 -0.019 0.03 0.019 ;
  LAYER v0 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m1 ;
    RECT -0.028 -0.021 0.028 0.021 ;
END V0_56x20_38H_56V

VIA V0_56x20_38H_70V
  LAYER m0 ;
    RECT -0.03 -0.019 0.03 0.019 ;
  LAYER v0 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m1 ;
    RECT -0.035 -0.021 0.035 0.021 ;
END V0_56x20_38H_70V

VIA V0_56x20_56H_35H
  LAYER m0 ;
    RECT -0.03 -0.028 0.03 0.028 ;
  LAYER v0 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m1 ;
    RECT -0.039 -0.0175 0.039 0.0175 ;
END V0_56x20_56H_35H

VIA V0_56x20_56H_56H
  LAYER m0 ;
    RECT -0.03 -0.028 0.03 0.028 ;
  LAYER v0 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m1 ;
    RECT -0.039 -0.028 0.039 0.028 ;
END V0_56x20_56H_56H

VIA V0_56x20_56H_56V
  LAYER m0 ;
    RECT -0.03 -0.028 0.03 0.028 ;
  LAYER v0 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m1 ;
    RECT -0.028 -0.021 0.028 0.021 ;
END V0_56x20_56H_56V

VIA V0_56x20_56H_70V
  LAYER m0 ;
    RECT -0.03 -0.028 0.03 0.028 ;
  LAYER v0 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m1 ;
    RECT -0.035 -0.021 0.035 0.021 ;
END V0_56x20_56H_70V

VIA V10_120x40S_120H_120V
  LAYER m10 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V10_120x40S_120H_120V

VIA V10_120x40S_120V_120V
  LAYER m10 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V10_120x40S_120V_120V

VIA V10_120x40S_160H_120V
  LAYER m10 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V10_120x40S_160H_120V

VIA V10_120x40S_160V_120V
  LAYER m10 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V10_120x40S_160V_120V

VIA V10_120x40S_200H_120V
  LAYER m10 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V10_120x40S_200H_120V

VIA V10_120x40S_200V_120V
  LAYER m10 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V10_120x40S_200V_120V

VIA V10_120x40S_40H_120V
  LAYER m10 ;
    RECT -0.084 -0.02 0.084 0.02 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V10_120x40S_40H_120V

VIA V10_120x40S_60H_120V
  LAYER m10 ;
    RECT -0.084 -0.03 0.084 0.03 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V10_120x40S_60H_120V

VIA V10_120x40S_80H_120V
  LAYER m10 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V10_120x40S_80H_120V

VIA V10_120x40_120H_120H
  LAYER m10 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V10_120x40_120H_120H

VIA V10_120x40_120H_160H
  LAYER m10 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V10_120x40_120H_160H

VIA V10_120x40_120H_160V
  LAYER m10 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V10_120x40_120H_160V

VIA V10_120x40_120H_200H
  LAYER m10 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V10_120x40_120H_200H

VIA V10_120x40_120H_200V
  LAYER m10 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V10_120x40_120H_200V

VIA V10_120x40_120H_240H
  LAYER m10 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.12 0.098 0.12 ;
END V10_120x40_120H_240H

VIA V10_120x40_120H_240V
  LAYER m10 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V10_120x40_120H_240V

VIA V10_120x40_160H_120H
  LAYER m10 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V10_120x40_160H_120H

VIA V10_120x40_160H_160H
  LAYER m10 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V10_120x40_160H_160H

VIA V10_120x40_160H_160V
  LAYER m10 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V10_120x40_160H_160V

VIA V10_120x40_160H_200H
  LAYER m10 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V10_120x40_160H_200H

VIA V10_120x40_160H_200V
  LAYER m10 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V10_120x40_160H_200V

VIA V10_120x40_160H_240H
  LAYER m10 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.12 0.098 0.12 ;
END V10_120x40_160H_240H

VIA V10_120x40_160H_240V
  LAYER m10 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V10_120x40_160H_240V

VIA V10_120x40_160V_120H
  LAYER m10 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V10_120x40_160V_120H

VIA V10_120x40_160V_160H
  LAYER m10 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V10_120x40_160V_160H

VIA V10_120x40_160V_160V
  LAYER m10 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V10_120x40_160V_160V

VIA V10_120x40_160V_200H
  LAYER m10 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V10_120x40_160V_200H

VIA V10_120x40_160V_200V
  LAYER m10 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V10_120x40_160V_200V

VIA V10_120x40_160V_240H
  LAYER m10 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.12 0.098 0.12 ;
END V10_120x40_160V_240H

VIA V10_120x40_160V_240V
  LAYER m10 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V10_120x40_160V_240V

VIA V10_120x40_200H_120H
  LAYER m10 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V10_120x40_200H_120H

VIA V10_120x40_200H_160H
  LAYER m10 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V10_120x40_200H_160H

VIA V10_120x40_200H_160V
  LAYER m10 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V10_120x40_200H_160V

VIA V10_120x40_200H_200H
  LAYER m10 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V10_120x40_200H_200H

VIA V10_120x40_200H_200V
  LAYER m10 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V10_120x40_200H_200V

VIA V10_120x40_200H_240H
  LAYER m10 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.12 0.098 0.12 ;
END V10_120x40_200H_240H

VIA V10_120x40_200H_240V
  LAYER m10 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V10_120x40_200H_240V

VIA V10_120x40_200V_120H
  LAYER m10 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V10_120x40_200V_120H

VIA V10_120x40_200V_160H
  LAYER m10 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V10_120x40_200V_160H

VIA V10_120x40_200V_160V
  LAYER m10 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V10_120x40_200V_160V

VIA V10_120x40_200V_200H
  LAYER m10 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V10_120x40_200V_200H

VIA V10_120x40_200V_200V
  LAYER m10 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V10_120x40_200V_200V

VIA V10_120x40_200V_240H
  LAYER m10 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.12 0.098 0.12 ;
END V10_120x40_200V_240H

VIA V10_120x40_200V_240V
  LAYER m10 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V10_120x40_200V_240V

VIA V10_120x40_80H_120H
  LAYER m10 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V10_120x40_80H_120H

VIA V10_120x40_80H_160H
  LAYER m10 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V10_120x40_80H_160H

VIA V10_120x40_80H_160V
  LAYER m10 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V10_120x40_80H_160V

VIA V10_120x40_80H_200H
  LAYER m10 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V10_120x40_80H_200H

VIA V10_120x40_80H_200V
  LAYER m10 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V10_120x40_80H_200V

VIA V10_120x40_80H_240H
  LAYER m10 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.098 -0.12 0.098 0.12 ;
END V10_120x40_80H_240H

VIA V10_120x40_80H_240V
  LAYER m10 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v10 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m11 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V10_120x40_80H_240V

VIA V10_120x60S_120H_120V
  LAYER m10 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v10 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m11 ;
    RECT -0.06 -0.068 0.06 0.068 ;
END V10_120x60S_120H_120V

VIA V10_120x60S_120V_120V
  LAYER m10 ;
    RECT -0.06 -0.054 0.06 0.054 ;
  LAYER v10 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m11 ;
    RECT -0.06 -0.068 0.06 0.068 ;
END V10_120x60S_120V_120V

VIA V10_120x60S_160H_120V
  LAYER m10 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v10 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m11 ;
    RECT -0.06 -0.068 0.06 0.068 ;
END V10_120x60S_160H_120V

VIA V10_120x60S_160V_120V
  LAYER m10 ;
    RECT -0.08 -0.054 0.08 0.054 ;
  LAYER v10 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m11 ;
    RECT -0.06 -0.068 0.06 0.068 ;
END V10_120x60S_160V_120V

VIA V10_120x60S_200H_120V
  LAYER m10 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v10 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m11 ;
    RECT -0.06 -0.068 0.06 0.068 ;
END V10_120x60S_200H_120V

VIA V10_120x60S_200V_120V
  LAYER m10 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v10 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m11 ;
    RECT -0.06 -0.068 0.06 0.068 ;
END V10_120x60S_200V_120V

VIA V10_120x60S_60H_120V
  LAYER m10 ;
    RECT -0.084 -0.03 0.084 0.03 ;
  LAYER v10 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m11 ;
    RECT -0.06 -0.068 0.06 0.068 ;
END V10_120x60S_60H_120V

VIA V10_120x60S_80H_120V
  LAYER m10 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v10 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m11 ;
    RECT -0.06 -0.068 0.06 0.068 ;
END V10_120x60S_80H_120V

VIA V10_160x40S_120H_160V
  LAYER m10 ;
    RECT -0.104 -0.06 0.104 0.06 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V10_160x40S_120H_160V

VIA V10_160x40S_160H_160V
  LAYER m10 ;
    RECT -0.104 -0.08 0.104 0.08 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V10_160x40S_160H_160V

VIA V10_160x40S_160V_160V
  LAYER m10 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V10_160x40S_160V_160V

VIA V10_160x40S_200H_160V
  LAYER m10 ;
    RECT -0.104 -0.1 0.104 0.1 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V10_160x40S_200H_160V

VIA V10_160x40S_200V_160V
  LAYER m10 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V10_160x40S_200V_160V

VIA V10_160x40S_40H_160V
  LAYER m10 ;
    RECT -0.104 -0.02 0.104 0.02 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V10_160x40S_40H_160V

VIA V10_160x40S_60H_160V
  LAYER m10 ;
    RECT -0.104 -0.03 0.104 0.03 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V10_160x40S_60H_160V

VIA V10_160x40S_80H_160V
  LAYER m10 ;
    RECT -0.104 -0.04 0.104 0.04 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V10_160x40S_80H_160V

VIA V10_160x40_120H_120H
  LAYER m10 ;
    RECT -0.104 -0.06 0.104 0.06 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.06 0.118 0.06 ;
END V10_160x40_120H_120H

VIA V10_160x40_120H_160H
  LAYER m10 ;
    RECT -0.104 -0.06 0.104 0.06 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.08 0.118 0.08 ;
END V10_160x40_120H_160H

VIA V10_160x40_120H_200H
  LAYER m10 ;
    RECT -0.104 -0.06 0.104 0.06 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.1 0.118 0.1 ;
END V10_160x40_120H_200H

VIA V10_160x40_120H_200V
  LAYER m10 ;
    RECT -0.104 -0.06 0.104 0.06 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V10_160x40_120H_200V

VIA V10_160x40_120H_240H
  LAYER m10 ;
    RECT -0.104 -0.06 0.104 0.06 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.12 0.118 0.12 ;
END V10_160x40_120H_240H

VIA V10_160x40_120H_240V
  LAYER m10 ;
    RECT -0.104 -0.06 0.104 0.06 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V10_160x40_120H_240V

VIA V10_160x40_160H_120H
  LAYER m10 ;
    RECT -0.104 -0.08 0.104 0.08 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.06 0.118 0.06 ;
END V10_160x40_160H_120H

VIA V10_160x40_160H_160H
  LAYER m10 ;
    RECT -0.104 -0.08 0.104 0.08 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.08 0.118 0.08 ;
END V10_160x40_160H_160H

VIA V10_160x40_160H_200H
  LAYER m10 ;
    RECT -0.104 -0.08 0.104 0.08 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.1 0.118 0.1 ;
END V10_160x40_160H_200H

VIA V10_160x40_160H_200V
  LAYER m10 ;
    RECT -0.104 -0.08 0.104 0.08 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V10_160x40_160H_200V

VIA V10_160x40_160H_240H
  LAYER m10 ;
    RECT -0.104 -0.08 0.104 0.08 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.12 0.118 0.12 ;
END V10_160x40_160H_240H

VIA V10_160x40_160H_240V
  LAYER m10 ;
    RECT -0.104 -0.08 0.104 0.08 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V10_160x40_160H_240V

VIA V10_160x40_200H_120H
  LAYER m10 ;
    RECT -0.104 -0.1 0.104 0.1 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.06 0.118 0.06 ;
END V10_160x40_200H_120H

VIA V10_160x40_200H_160H
  LAYER m10 ;
    RECT -0.104 -0.1 0.104 0.1 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.08 0.118 0.08 ;
END V10_160x40_200H_160H

VIA V10_160x40_200H_200H
  LAYER m10 ;
    RECT -0.104 -0.1 0.104 0.1 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.1 0.118 0.1 ;
END V10_160x40_200H_200H

VIA V10_160x40_200H_200V
  LAYER m10 ;
    RECT -0.104 -0.1 0.104 0.1 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V10_160x40_200H_200V

VIA V10_160x40_200H_240H
  LAYER m10 ;
    RECT -0.104 -0.1 0.104 0.1 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.12 0.118 0.12 ;
END V10_160x40_200H_240H

VIA V10_160x40_200H_240V
  LAYER m10 ;
    RECT -0.104 -0.1 0.104 0.1 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V10_160x40_200H_240V

VIA V10_160x40_200V_120H
  LAYER m10 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.06 0.118 0.06 ;
END V10_160x40_200V_120H

VIA V10_160x40_200V_160H
  LAYER m10 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.08 0.118 0.08 ;
END V10_160x40_200V_160H

VIA V10_160x40_200V_200H
  LAYER m10 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.1 0.118 0.1 ;
END V10_160x40_200V_200H

VIA V10_160x40_200V_200V
  LAYER m10 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V10_160x40_200V_200V

VIA V10_160x40_200V_240H
  LAYER m10 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.12 0.118 0.12 ;
END V10_160x40_200V_240H

VIA V10_160x40_200V_240V
  LAYER m10 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V10_160x40_200V_240V

VIA V10_160x40_80H_120H
  LAYER m10 ;
    RECT -0.104 -0.04 0.104 0.04 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.06 0.118 0.06 ;
END V10_160x40_80H_120H

VIA V10_160x40_80H_160H
  LAYER m10 ;
    RECT -0.104 -0.04 0.104 0.04 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.08 0.118 0.08 ;
END V10_160x40_80H_160H

VIA V10_160x40_80H_200H
  LAYER m10 ;
    RECT -0.104 -0.04 0.104 0.04 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.1 0.118 0.1 ;
END V10_160x40_80H_200H

VIA V10_160x40_80H_200V
  LAYER m10 ;
    RECT -0.104 -0.04 0.104 0.04 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V10_160x40_80H_200V

VIA V10_160x40_80H_240H
  LAYER m10 ;
    RECT -0.104 -0.04 0.104 0.04 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.118 -0.12 0.118 0.12 ;
END V10_160x40_80H_240H

VIA V10_160x40_80H_240V
  LAYER m10 ;
    RECT -0.104 -0.04 0.104 0.04 ;
  LAYER v10 ;
    RECT -0.08 -0.02 0.08 0.02 ;
  LAYER m11 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V10_160x40_80H_240V

VIA V10_40Sx120_120H_120H
  LAYER m10 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V10_40Sx120_120H_120H

VIA V10_40Sx120_120V_120H
  LAYER m10 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V10_40Sx120_120V_120H

VIA V10_40Sx120_160H_120H
  LAYER m10 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V10_40Sx120_160H_120H

VIA V10_40Sx120_160V_120H
  LAYER m10 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V10_40Sx120_160V_120H

VIA V10_40Sx120_200H_120H
  LAYER m10 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V10_40Sx120_200H_120H

VIA V10_40Sx120_200V_120H
  LAYER m10 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V10_40Sx120_200V_120H

VIA V10_40Sx120_80V_120H
  LAYER m10 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V10_40Sx120_80V_120H

VIA V10_40x120_120V_120V
  LAYER m10 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V10_40x120_120V_120V

VIA V10_40x120_120V_160H
  LAYER m10 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V10_40x120_120V_160H

VIA V10_40x120_120V_160V
  LAYER m10 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V10_40x120_120V_160V

VIA V10_40x120_120V_200H
  LAYER m10 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V10_40x120_120V_200H

VIA V10_40x120_120V_200V
  LAYER m10 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V10_40x120_120V_200V

VIA V10_40x120_120V_240H
  LAYER m10 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V10_40x120_120V_240H

VIA V10_40x120_120V_240V
  LAYER m10 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.12 -0.098 0.12 0.098 ;
END V10_40x120_120V_240V

VIA V10_40x120_120V_90V
  LAYER m10 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.045 -0.098 0.045 0.098 ;
END V10_40x120_120V_90V

VIA V10_40x120_160H_120V
  LAYER m10 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V10_40x120_160H_120V

VIA V10_40x120_160H_160H
  LAYER m10 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V10_40x120_160H_160H

VIA V10_40x120_160H_160V
  LAYER m10 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V10_40x120_160H_160V

VIA V10_40x120_160H_200H
  LAYER m10 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V10_40x120_160H_200H

VIA V10_40x120_160H_200V
  LAYER m10 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V10_40x120_160H_200V

VIA V10_40x120_160H_240H
  LAYER m10 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V10_40x120_160H_240H

VIA V10_40x120_160H_240V
  LAYER m10 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.12 -0.098 0.12 0.098 ;
END V10_40x120_160H_240V

VIA V10_40x120_160H_90V
  LAYER m10 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.045 -0.098 0.045 0.098 ;
END V10_40x120_160H_90V

VIA V10_40x120_160V_120V
  LAYER m10 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V10_40x120_160V_120V

VIA V10_40x120_160V_160H
  LAYER m10 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V10_40x120_160V_160H

VIA V10_40x120_160V_160V
  LAYER m10 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V10_40x120_160V_160V

VIA V10_40x120_160V_200H
  LAYER m10 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V10_40x120_160V_200H

VIA V10_40x120_160V_200V
  LAYER m10 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V10_40x120_160V_200V

VIA V10_40x120_160V_240H
  LAYER m10 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V10_40x120_160V_240H

VIA V10_40x120_160V_240V
  LAYER m10 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.12 -0.098 0.12 0.098 ;
END V10_40x120_160V_240V

VIA V10_40x120_160V_90V
  LAYER m10 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.045 -0.098 0.045 0.098 ;
END V10_40x120_160V_90V

VIA V10_40x120_200H_120V
  LAYER m10 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V10_40x120_200H_120V

VIA V10_40x120_200H_160H
  LAYER m10 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V10_40x120_200H_160H

VIA V10_40x120_200H_160V
  LAYER m10 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V10_40x120_200H_160V

VIA V10_40x120_200H_200H
  LAYER m10 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V10_40x120_200H_200H

VIA V10_40x120_200H_200V
  LAYER m10 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V10_40x120_200H_200V

VIA V10_40x120_200H_240H
  LAYER m10 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V10_40x120_200H_240H

VIA V10_40x120_200H_240V
  LAYER m10 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.12 -0.098 0.12 0.098 ;
END V10_40x120_200H_240V

VIA V10_40x120_200H_90V
  LAYER m10 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.045 -0.098 0.045 0.098 ;
END V10_40x120_200H_90V

VIA V10_40x120_200V_120V
  LAYER m10 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V10_40x120_200V_120V

VIA V10_40x120_200V_160H
  LAYER m10 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V10_40x120_200V_160H

VIA V10_40x120_200V_160V
  LAYER m10 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V10_40x120_200V_160V

VIA V10_40x120_200V_200H
  LAYER m10 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V10_40x120_200V_200H

VIA V10_40x120_200V_200V
  LAYER m10 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V10_40x120_200V_200V

VIA V10_40x120_200V_240H
  LAYER m10 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V10_40x120_200V_240H

VIA V10_40x120_200V_240V
  LAYER m10 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.12 -0.098 0.12 0.098 ;
END V10_40x120_200V_240V

VIA V10_40x120_200V_90V
  LAYER m10 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.045 -0.098 0.045 0.098 ;
END V10_40x120_200V_90V

VIA V10_40x120_80V_120V
  LAYER m10 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V10_40x120_80V_120V

VIA V10_40x120_80V_160H
  LAYER m10 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V10_40x120_80V_160H

VIA V10_40x120_80V_160V
  LAYER m10 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V10_40x120_80V_160V

VIA V10_40x120_80V_200H
  LAYER m10 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V10_40x120_80V_200H

VIA V10_40x120_80V_200V
  LAYER m10 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V10_40x120_80V_200V

VIA V10_40x120_80V_240H
  LAYER m10 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V10_40x120_80V_240H

VIA V10_40x120_80V_240V
  LAYER m10 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.12 -0.098 0.12 0.098 ;
END V10_40x120_80V_240V

VIA V10_40x120_80V_90V
  LAYER m10 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v10 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m11 ;
    RECT -0.045 -0.098 0.045 0.098 ;
END V10_40x120_80V_90V

VIA V10_40x160_120V_120V
  LAYER m10 ;
    RECT -0.06 -0.104 0.06 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.06 -0.118 0.06 0.118 ;
END V10_40x160_120V_120V

VIA V10_40x160_120V_160V
  LAYER m10 ;
    RECT -0.06 -0.104 0.06 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.08 -0.118 0.08 0.118 ;
END V10_40x160_120V_160V

VIA V10_40x160_120V_200H
  LAYER m10 ;
    RECT -0.06 -0.104 0.06 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V10_40x160_120V_200H

VIA V10_40x160_120V_200V
  LAYER m10 ;
    RECT -0.06 -0.104 0.06 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.1 -0.118 0.1 0.118 ;
END V10_40x160_120V_200V

VIA V10_40x160_120V_240H
  LAYER m10 ;
    RECT -0.06 -0.104 0.06 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V10_40x160_120V_240H

VIA V10_40x160_120V_240V
  LAYER m10 ;
    RECT -0.06 -0.104 0.06 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.12 -0.118 0.12 0.118 ;
END V10_40x160_120V_240V

VIA V10_40x160_120V_90V
  LAYER m10 ;
    RECT -0.06 -0.104 0.06 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.045 -0.118 0.045 0.118 ;
END V10_40x160_120V_90V

VIA V10_40x160_160V_120V
  LAYER m10 ;
    RECT -0.08 -0.104 0.08 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.06 -0.118 0.06 0.118 ;
END V10_40x160_160V_120V

VIA V10_40x160_160V_160V
  LAYER m10 ;
    RECT -0.08 -0.104 0.08 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.08 -0.118 0.08 0.118 ;
END V10_40x160_160V_160V

VIA V10_40x160_160V_200H
  LAYER m10 ;
    RECT -0.08 -0.104 0.08 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V10_40x160_160V_200H

VIA V10_40x160_160V_200V
  LAYER m10 ;
    RECT -0.08 -0.104 0.08 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.1 -0.118 0.1 0.118 ;
END V10_40x160_160V_200V

VIA V10_40x160_160V_240H
  LAYER m10 ;
    RECT -0.08 -0.104 0.08 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V10_40x160_160V_240H

VIA V10_40x160_160V_240V
  LAYER m10 ;
    RECT -0.08 -0.104 0.08 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.12 -0.118 0.12 0.118 ;
END V10_40x160_160V_240V

VIA V10_40x160_160V_90V
  LAYER m10 ;
    RECT -0.08 -0.104 0.08 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.045 -0.118 0.045 0.118 ;
END V10_40x160_160V_90V

VIA V10_40x160_200H_120V
  LAYER m10 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.06 -0.118 0.06 0.118 ;
END V10_40x160_200H_120V

VIA V10_40x160_200H_160V
  LAYER m10 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.08 -0.118 0.08 0.118 ;
END V10_40x160_200H_160V

VIA V10_40x160_200H_200H
  LAYER m10 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V10_40x160_200H_200H

VIA V10_40x160_200H_200V
  LAYER m10 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.1 -0.118 0.1 0.118 ;
END V10_40x160_200H_200V

VIA V10_40x160_200H_240H
  LAYER m10 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V10_40x160_200H_240H

VIA V10_40x160_200H_240V
  LAYER m10 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.12 -0.118 0.12 0.118 ;
END V10_40x160_200H_240V

VIA V10_40x160_200H_90V
  LAYER m10 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.045 -0.118 0.045 0.118 ;
END V10_40x160_200H_90V

VIA V10_40x160_200V_120V
  LAYER m10 ;
    RECT -0.1 -0.104 0.1 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.06 -0.118 0.06 0.118 ;
END V10_40x160_200V_120V

VIA V10_40x160_200V_160V
  LAYER m10 ;
    RECT -0.1 -0.104 0.1 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.08 -0.118 0.08 0.118 ;
END V10_40x160_200V_160V

VIA V10_40x160_200V_200H
  LAYER m10 ;
    RECT -0.1 -0.104 0.1 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V10_40x160_200V_200H

VIA V10_40x160_200V_200V
  LAYER m10 ;
    RECT -0.1 -0.104 0.1 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.1 -0.118 0.1 0.118 ;
END V10_40x160_200V_200V

VIA V10_40x160_200V_240H
  LAYER m10 ;
    RECT -0.1 -0.104 0.1 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V10_40x160_200V_240H

VIA V10_40x160_200V_240V
  LAYER m10 ;
    RECT -0.1 -0.104 0.1 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.12 -0.118 0.12 0.118 ;
END V10_40x160_200V_240V

VIA V10_40x160_200V_90V
  LAYER m10 ;
    RECT -0.1 -0.104 0.1 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.045 -0.118 0.045 0.118 ;
END V10_40x160_200V_90V

VIA V10_40x160_80V_120V
  LAYER m10 ;
    RECT -0.04 -0.104 0.04 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.06 -0.118 0.06 0.118 ;
END V10_40x160_80V_120V

VIA V10_40x160_80V_160V
  LAYER m10 ;
    RECT -0.04 -0.104 0.04 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.08 -0.118 0.08 0.118 ;
END V10_40x160_80V_160V

VIA V10_40x160_80V_200H
  LAYER m10 ;
    RECT -0.04 -0.104 0.04 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V10_40x160_80V_200H

VIA V10_40x160_80V_200V
  LAYER m10 ;
    RECT -0.04 -0.104 0.04 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.1 -0.118 0.1 0.118 ;
END V10_40x160_80V_200V

VIA V10_40x160_80V_240H
  LAYER m10 ;
    RECT -0.04 -0.104 0.04 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V10_40x160_80V_240H

VIA V10_40x160_80V_240V
  LAYER m10 ;
    RECT -0.04 -0.104 0.04 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.12 -0.118 0.12 0.118 ;
END V10_40x160_80V_240V

VIA V10_40x160_80V_90V
  LAYER m10 ;
    RECT -0.04 -0.104 0.04 0.104 ;
  LAYER v10 ;
    RECT -0.02 -0.08 0.02 0.08 ;
  LAYER m11 ;
    RECT -0.045 -0.118 0.045 0.118 ;
END V10_40x160_80V_90V

VIA V10_60x40S_120H_60V
  LAYER m10 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v10 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m11 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V10_60x40S_120H_60V

VIA V10_60x40S_120V_60V
  LAYER m10 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v10 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m11 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V10_60x40S_120V_60V

VIA V10_60x40S_160H_60V
  LAYER m10 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v10 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m11 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V10_60x40S_160H_60V

VIA V10_60x40S_160V_60V
  LAYER m10 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v10 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m11 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V10_60x40S_160V_60V

VIA V10_60x40S_200H_60V
  LAYER m10 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v10 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m11 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V10_60x40S_200H_60V

VIA V10_60x40S_200V_60V
  LAYER m10 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v10 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m11 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V10_60x40S_200V_60V

VIA V10_60x40S_40H_60V
  LAYER m10 ;
    RECT -0.054 -0.02 0.054 0.02 ;
  LAYER v10 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m11 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V10_60x40S_40H_60V

VIA V10_60x40S_60H_60V
  LAYER m10 ;
    RECT -0.054 -0.03 0.054 0.03 ;
  LAYER v10 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m11 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V10_60x40S_60H_60V

VIA V10_60x40S_80H_60V
  LAYER m10 ;
    RECT -0.054 -0.04 0.054 0.04 ;
  LAYER v10 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m11 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V10_60x40S_80H_60V

VIA V10_60x40S_80V_60V
  LAYER m10 ;
    RECT -0.04 -0.044 0.04 0.044 ;
  LAYER v10 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m11 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V10_60x40S_80V_60V

VIA V10_60x60S_120H_60V
  LAYER m10 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v10 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m11 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V10_60x60S_120H_60V

VIA V10_60x60S_120V_60V
  LAYER m10 ;
    RECT -0.06 -0.054 0.06 0.054 ;
  LAYER v10 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m11 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V10_60x60S_120V_60V

VIA V10_60x60S_160H_60V
  LAYER m10 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v10 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m11 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V10_60x60S_160H_60V

VIA V10_60x60S_160V_60V
  LAYER m10 ;
    RECT -0.08 -0.054 0.08 0.054 ;
  LAYER v10 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m11 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V10_60x60S_160V_60V

VIA V10_60x60S_200H_60V
  LAYER m10 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v10 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m11 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V10_60x60S_200H_60V

VIA V10_60x60S_200V_60V
  LAYER m10 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v10 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m11 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V10_60x60S_200V_60V

VIA V10_60x60S_60H_60V
  LAYER m10 ;
    RECT -0.054 -0.03 0.054 0.03 ;
  LAYER v10 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m11 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V10_60x60S_60H_60V

VIA V10_60x60S_80H_60V
  LAYER m10 ;
    RECT -0.054 -0.04 0.054 0.04 ;
  LAYER v10 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m11 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V10_60x60S_80H_60V

VIA V10_60x60S_80V_60V
  LAYER m10 ;
    RECT -0.04 -0.054 0.04 0.054 ;
  LAYER v10 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m11 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V10_60x60S_80V_60V

VIA V10_90x40S_120H_90V
  LAYER m10 ;
    RECT -0.069 -0.06 0.069 0.06 ;
  LAYER v10 ;
    RECT -0.045 -0.02 0.045 0.02 ;
  LAYER m11 ;
    RECT -0.045 -0.058 0.045 0.058 ;
END V10_90x40S_120H_90V

VIA V10_90x40S_120V_90V
  LAYER m10 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v10 ;
    RECT -0.045 -0.02 0.045 0.02 ;
  LAYER m11 ;
    RECT -0.045 -0.058 0.045 0.058 ;
END V10_90x40S_120V_90V

VIA V10_90x40S_160H_90V
  LAYER m10 ;
    RECT -0.069 -0.08 0.069 0.08 ;
  LAYER v10 ;
    RECT -0.045 -0.02 0.045 0.02 ;
  LAYER m11 ;
    RECT -0.045 -0.058 0.045 0.058 ;
END V10_90x40S_160H_90V

VIA V10_90x40S_160V_90V
  LAYER m10 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v10 ;
    RECT -0.045 -0.02 0.045 0.02 ;
  LAYER m11 ;
    RECT -0.045 -0.058 0.045 0.058 ;
END V10_90x40S_160V_90V

VIA V10_90x40S_200H_90V
  LAYER m10 ;
    RECT -0.069 -0.1 0.069 0.1 ;
  LAYER v10 ;
    RECT -0.045 -0.02 0.045 0.02 ;
  LAYER m11 ;
    RECT -0.045 -0.058 0.045 0.058 ;
END V10_90x40S_200H_90V

VIA V10_90x40S_200V_90V
  LAYER m10 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v10 ;
    RECT -0.045 -0.02 0.045 0.02 ;
  LAYER m11 ;
    RECT -0.045 -0.058 0.045 0.058 ;
END V10_90x40S_200V_90V

VIA V10_90x40S_40H_90V
  LAYER m10 ;
    RECT -0.069 -0.02 0.069 0.02 ;
  LAYER v10 ;
    RECT -0.045 -0.02 0.045 0.02 ;
  LAYER m11 ;
    RECT -0.045 -0.058 0.045 0.058 ;
END V10_90x40S_40H_90V

VIA V10_90x40S_60H_90V
  LAYER m10 ;
    RECT -0.069 -0.03 0.069 0.03 ;
  LAYER v10 ;
    RECT -0.045 -0.02 0.045 0.02 ;
  LAYER m11 ;
    RECT -0.045 -0.058 0.045 0.058 ;
END V10_90x40S_60H_90V

VIA V10_90x40S_80H_90V
  LAYER m10 ;
    RECT -0.069 -0.04 0.069 0.04 ;
  LAYER v10 ;
    RECT -0.045 -0.02 0.045 0.02 ;
  LAYER m11 ;
    RECT -0.045 -0.058 0.045 0.058 ;
END V10_90x40S_80H_90V

VIA V10_90x60S_120H_90V
  LAYER m10 ;
    RECT -0.069 -0.06 0.069 0.06 ;
  LAYER v10 ;
    RECT -0.045 -0.03 0.045 0.03 ;
  LAYER m11 ;
    RECT -0.045 -0.068 0.045 0.068 ;
END V10_90x60S_120H_90V

VIA V10_90x60S_120V_90V
  LAYER m10 ;
    RECT -0.06 -0.054 0.06 0.054 ;
  LAYER v10 ;
    RECT -0.045 -0.03 0.045 0.03 ;
  LAYER m11 ;
    RECT -0.045 -0.068 0.045 0.068 ;
END V10_90x60S_120V_90V

VIA V10_90x60S_160H_90V
  LAYER m10 ;
    RECT -0.069 -0.08 0.069 0.08 ;
  LAYER v10 ;
    RECT -0.045 -0.03 0.045 0.03 ;
  LAYER m11 ;
    RECT -0.045 -0.068 0.045 0.068 ;
END V10_90x60S_160H_90V

VIA V10_90x60S_160V_90V
  LAYER m10 ;
    RECT -0.08 -0.054 0.08 0.054 ;
  LAYER v10 ;
    RECT -0.045 -0.03 0.045 0.03 ;
  LAYER m11 ;
    RECT -0.045 -0.068 0.045 0.068 ;
END V10_90x60S_160V_90V

VIA V10_90x60S_200H_90V
  LAYER m10 ;
    RECT -0.069 -0.1 0.069 0.1 ;
  LAYER v10 ;
    RECT -0.045 -0.03 0.045 0.03 ;
  LAYER m11 ;
    RECT -0.045 -0.068 0.045 0.068 ;
END V10_90x60S_200H_90V

VIA V10_90x60S_200V_90V
  LAYER m10 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v10 ;
    RECT -0.045 -0.03 0.045 0.03 ;
  LAYER m11 ;
    RECT -0.045 -0.068 0.045 0.068 ;
END V10_90x60S_200V_90V

VIA V10_90x60S_60H_90V
  LAYER m10 ;
    RECT -0.069 -0.03 0.069 0.03 ;
  LAYER v10 ;
    RECT -0.045 -0.03 0.045 0.03 ;
  LAYER m11 ;
    RECT -0.045 -0.068 0.045 0.068 ;
END V10_90x60S_60H_90V

VIA V10_90x60S_80H_90V
  LAYER m10 ;
    RECT -0.069 -0.04 0.069 0.04 ;
  LAYER v10 ;
    RECT -0.045 -0.03 0.045 0.03 ;
  LAYER m11 ;
    RECT -0.045 -0.068 0.045 0.068 ;
END V10_90x60S_80H_90V

VIA V11_120x40S_120H_120V
  LAYER m11 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V11_120x40S_120H_120V

VIA V11_120x40S_120V_120V
  LAYER m11 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V11_120x40S_120V_120V

VIA V11_120x40S_160H_120V
  LAYER m11 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V11_120x40S_160H_120V

VIA V11_120x40S_160V_120V
  LAYER m11 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V11_120x40S_160V_120V

VIA V11_120x40S_200H_120V
  LAYER m11 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V11_120x40S_200H_120V

VIA V11_120x40S_200V_120V
  LAYER m11 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V11_120x40S_200V_120V

VIA V11_120x40S_240H_120V
  LAYER m11 ;
    RECT -0.084 -0.12 0.084 0.12 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V11_120x40S_240H_120V

VIA V11_120x40S_240V_120V
  LAYER m11 ;
    RECT -0.12 -0.044 0.12 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V11_120x40S_240V_120V

VIA V11_120x40_120H_120H
  LAYER m11 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V11_120x40_120H_120H

VIA V11_120x40_120H_160H
  LAYER m11 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V11_120x40_120H_160H

VIA V11_120x40_120H_160V
  LAYER m11 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V11_120x40_120H_160V

VIA V11_120x40_120H_200H
  LAYER m11 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V11_120x40_120H_200H

VIA V11_120x40_120H_200V
  LAYER m11 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V11_120x40_120H_200V

VIA V11_120x40_120H_240H
  LAYER m11 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.12 0.098 0.12 ;
END V11_120x40_120H_240H

VIA V11_120x40_120H_240V
  LAYER m11 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V11_120x40_120H_240V

VIA V11_120x40_120H_90H
  LAYER m11 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.045 0.098 0.045 ;
END V11_120x40_120H_90H

VIA V11_120x40_160H_120H
  LAYER m11 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V11_120x40_160H_120H

VIA V11_120x40_160H_160H
  LAYER m11 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V11_120x40_160H_160H

VIA V11_120x40_160H_160V
  LAYER m11 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V11_120x40_160H_160V

VIA V11_120x40_160H_200H
  LAYER m11 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V11_120x40_160H_200H

VIA V11_120x40_160H_200V
  LAYER m11 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V11_120x40_160H_200V

VIA V11_120x40_160H_240H
  LAYER m11 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.12 0.098 0.12 ;
END V11_120x40_160H_240H

VIA V11_120x40_160H_240V
  LAYER m11 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V11_120x40_160H_240V

VIA V11_120x40_160H_90H
  LAYER m11 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.045 0.098 0.045 ;
END V11_120x40_160H_90H

VIA V11_120x40_160V_120H
  LAYER m11 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V11_120x40_160V_120H

VIA V11_120x40_160V_160H
  LAYER m11 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V11_120x40_160V_160H

VIA V11_120x40_160V_160V
  LAYER m11 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V11_120x40_160V_160V

VIA V11_120x40_160V_200H
  LAYER m11 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V11_120x40_160V_200H

VIA V11_120x40_160V_200V
  LAYER m11 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V11_120x40_160V_200V

VIA V11_120x40_160V_240H
  LAYER m11 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.12 0.098 0.12 ;
END V11_120x40_160V_240H

VIA V11_120x40_160V_240V
  LAYER m11 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V11_120x40_160V_240V

VIA V11_120x40_160V_90H
  LAYER m11 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.045 0.098 0.045 ;
END V11_120x40_160V_90H

VIA V11_120x40_200H_120H
  LAYER m11 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V11_120x40_200H_120H

VIA V11_120x40_200H_160H
  LAYER m11 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V11_120x40_200H_160H

VIA V11_120x40_200H_160V
  LAYER m11 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V11_120x40_200H_160V

VIA V11_120x40_200H_200H
  LAYER m11 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V11_120x40_200H_200H

VIA V11_120x40_200H_200V
  LAYER m11 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V11_120x40_200H_200V

VIA V11_120x40_200H_240H
  LAYER m11 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.12 0.098 0.12 ;
END V11_120x40_200H_240H

VIA V11_120x40_200H_240V
  LAYER m11 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V11_120x40_200H_240V

VIA V11_120x40_200H_90H
  LAYER m11 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.045 0.098 0.045 ;
END V11_120x40_200H_90H

VIA V11_120x40_200V_120H
  LAYER m11 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V11_120x40_200V_120H

VIA V11_120x40_200V_160H
  LAYER m11 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V11_120x40_200V_160H

VIA V11_120x40_200V_160V
  LAYER m11 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V11_120x40_200V_160V

VIA V11_120x40_200V_200H
  LAYER m11 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V11_120x40_200V_200H

VIA V11_120x40_200V_200V
  LAYER m11 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V11_120x40_200V_200V

VIA V11_120x40_200V_240H
  LAYER m11 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.12 0.098 0.12 ;
END V11_120x40_200V_240H

VIA V11_120x40_200V_240V
  LAYER m11 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V11_120x40_200V_240V

VIA V11_120x40_200V_90H
  LAYER m11 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.045 0.098 0.045 ;
END V11_120x40_200V_90H

VIA V11_120x40_240H_120H
  LAYER m11 ;
    RECT -0.084 -0.12 0.084 0.12 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V11_120x40_240H_120H

VIA V11_120x40_240H_160H
  LAYER m11 ;
    RECT -0.084 -0.12 0.084 0.12 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V11_120x40_240H_160H

VIA V11_120x40_240H_160V
  LAYER m11 ;
    RECT -0.084 -0.12 0.084 0.12 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V11_120x40_240H_160V

VIA V11_120x40_240H_200H
  LAYER m11 ;
    RECT -0.084 -0.12 0.084 0.12 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V11_120x40_240H_200H

VIA V11_120x40_240H_200V
  LAYER m11 ;
    RECT -0.084 -0.12 0.084 0.12 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V11_120x40_240H_200V

VIA V11_120x40_240H_240H
  LAYER m11 ;
    RECT -0.084 -0.12 0.084 0.12 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.12 0.098 0.12 ;
END V11_120x40_240H_240H

VIA V11_120x40_240H_240V
  LAYER m11 ;
    RECT -0.084 -0.12 0.084 0.12 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V11_120x40_240H_240V

VIA V11_120x40_240H_90H
  LAYER m11 ;
    RECT -0.084 -0.12 0.084 0.12 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.045 0.098 0.045 ;
END V11_120x40_240H_90H

VIA V11_120x40_240V_120H
  LAYER m11 ;
    RECT -0.12 -0.044 0.12 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V11_120x40_240V_120H

VIA V11_120x40_240V_160H
  LAYER m11 ;
    RECT -0.12 -0.044 0.12 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V11_120x40_240V_160H

VIA V11_120x40_240V_160V
  LAYER m11 ;
    RECT -0.12 -0.044 0.12 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V11_120x40_240V_160V

VIA V11_120x40_240V_200H
  LAYER m11 ;
    RECT -0.12 -0.044 0.12 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V11_120x40_240V_200H

VIA V11_120x40_240V_200V
  LAYER m11 ;
    RECT -0.12 -0.044 0.12 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V11_120x40_240V_200V

VIA V11_120x40_240V_240H
  LAYER m11 ;
    RECT -0.12 -0.044 0.12 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.12 0.098 0.12 ;
END V11_120x40_240V_240H

VIA V11_120x40_240V_240V
  LAYER m11 ;
    RECT -0.12 -0.044 0.12 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.12 -0.058 0.12 0.058 ;
END V11_120x40_240V_240V

VIA V11_120x40_240V_90H
  LAYER m11 ;
    RECT -0.12 -0.044 0.12 0.044 ;
  LAYER v11 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m12 ;
    RECT -0.098 -0.045 0.098 0.045 ;
END V11_120x40_240V_90H

VIA V11_160x60_120H_120H
  LAYER m11 ;
    RECT -0.104 -0.06 0.104 0.06 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.06 0.118 0.06 ;
END V11_160x60_120H_120H

VIA V11_160x60_120H_160H
  LAYER m11 ;
    RECT -0.104 -0.06 0.104 0.06 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.08 0.118 0.08 ;
END V11_160x60_120H_160H

VIA V11_160x60_120H_200H
  LAYER m11 ;
    RECT -0.104 -0.06 0.104 0.06 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.1 0.118 0.1 ;
END V11_160x60_120H_200H

VIA V11_160x60_120H_200V
  LAYER m11 ;
    RECT -0.104 -0.06 0.104 0.06 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.1 -0.068 0.1 0.068 ;
END V11_160x60_120H_200V

VIA V11_160x60_120H_240H
  LAYER m11 ;
    RECT -0.104 -0.06 0.104 0.06 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.12 0.118 0.12 ;
END V11_160x60_120H_240H

VIA V11_160x60_120H_240V
  LAYER m11 ;
    RECT -0.104 -0.06 0.104 0.06 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.12 -0.068 0.12 0.068 ;
END V11_160x60_120H_240V

VIA V11_160x60_160H_120H
  LAYER m11 ;
    RECT -0.104 -0.08 0.104 0.08 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.06 0.118 0.06 ;
END V11_160x60_160H_120H

VIA V11_160x60_160H_160H
  LAYER m11 ;
    RECT -0.104 -0.08 0.104 0.08 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.08 0.118 0.08 ;
END V11_160x60_160H_160H

VIA V11_160x60_160H_200H
  LAYER m11 ;
    RECT -0.104 -0.08 0.104 0.08 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.1 0.118 0.1 ;
END V11_160x60_160H_200H

VIA V11_160x60_160H_200V
  LAYER m11 ;
    RECT -0.104 -0.08 0.104 0.08 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.1 -0.068 0.1 0.068 ;
END V11_160x60_160H_200V

VIA V11_160x60_160H_240H
  LAYER m11 ;
    RECT -0.104 -0.08 0.104 0.08 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.12 0.118 0.12 ;
END V11_160x60_160H_240H

VIA V11_160x60_160H_240V
  LAYER m11 ;
    RECT -0.104 -0.08 0.104 0.08 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.12 -0.068 0.12 0.068 ;
END V11_160x60_160H_240V

VIA V11_160x60_200H_120H
  LAYER m11 ;
    RECT -0.104 -0.1 0.104 0.1 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.06 0.118 0.06 ;
END V11_160x60_200H_120H

VIA V11_160x60_200H_160H
  LAYER m11 ;
    RECT -0.104 -0.1 0.104 0.1 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.08 0.118 0.08 ;
END V11_160x60_200H_160H

VIA V11_160x60_200H_200H
  LAYER m11 ;
    RECT -0.104 -0.1 0.104 0.1 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.1 0.118 0.1 ;
END V11_160x60_200H_200H

VIA V11_160x60_200H_200V
  LAYER m11 ;
    RECT -0.104 -0.1 0.104 0.1 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.1 -0.068 0.1 0.068 ;
END V11_160x60_200H_200V

VIA V11_160x60_200H_240H
  LAYER m11 ;
    RECT -0.104 -0.1 0.104 0.1 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.12 0.118 0.12 ;
END V11_160x60_200H_240H

VIA V11_160x60_200H_240V
  LAYER m11 ;
    RECT -0.104 -0.1 0.104 0.1 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.12 -0.068 0.12 0.068 ;
END V11_160x60_200H_240V

VIA V11_160x60_200V_120H
  LAYER m11 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.06 0.118 0.06 ;
END V11_160x60_200V_120H

VIA V11_160x60_200V_160H
  LAYER m11 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.08 0.118 0.08 ;
END V11_160x60_200V_160H

VIA V11_160x60_200V_200H
  LAYER m11 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.1 0.118 0.1 ;
END V11_160x60_200V_200H

VIA V11_160x60_200V_200V
  LAYER m11 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.1 -0.068 0.1 0.068 ;
END V11_160x60_200V_200V

VIA V11_160x60_200V_240H
  LAYER m11 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.12 0.118 0.12 ;
END V11_160x60_200V_240H

VIA V11_160x60_200V_240V
  LAYER m11 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.12 -0.068 0.12 0.068 ;
END V11_160x60_200V_240V

VIA V11_160x60_240H_120H
  LAYER m11 ;
    RECT -0.104 -0.12 0.104 0.12 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.06 0.118 0.06 ;
END V11_160x60_240H_120H

VIA V11_160x60_240H_160H
  LAYER m11 ;
    RECT -0.104 -0.12 0.104 0.12 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.08 0.118 0.08 ;
END V11_160x60_240H_160H

VIA V11_160x60_240H_200H
  LAYER m11 ;
    RECT -0.104 -0.12 0.104 0.12 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.1 0.118 0.1 ;
END V11_160x60_240H_200H

VIA V11_160x60_240H_200V
  LAYER m11 ;
    RECT -0.104 -0.12 0.104 0.12 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.1 -0.068 0.1 0.068 ;
END V11_160x60_240H_200V

VIA V11_160x60_240H_240H
  LAYER m11 ;
    RECT -0.104 -0.12 0.104 0.12 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.12 0.118 0.12 ;
END V11_160x60_240H_240H

VIA V11_160x60_240H_240V
  LAYER m11 ;
    RECT -0.104 -0.12 0.104 0.12 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.12 -0.068 0.12 0.068 ;
END V11_160x60_240H_240V

VIA V11_160x60_240V_120H
  LAYER m11 ;
    RECT -0.12 -0.054 0.12 0.054 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.06 0.118 0.06 ;
END V11_160x60_240V_120H

VIA V11_160x60_240V_160H
  LAYER m11 ;
    RECT -0.12 -0.054 0.12 0.054 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.08 0.118 0.08 ;
END V11_160x60_240V_160H

VIA V11_160x60_240V_200H
  LAYER m11 ;
    RECT -0.12 -0.054 0.12 0.054 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.1 0.118 0.1 ;
END V11_160x60_240V_200H

VIA V11_160x60_240V_200V
  LAYER m11 ;
    RECT -0.12 -0.054 0.12 0.054 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.1 -0.068 0.1 0.068 ;
END V11_160x60_240V_200V

VIA V11_160x60_240V_240H
  LAYER m11 ;
    RECT -0.12 -0.054 0.12 0.054 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.118 -0.12 0.118 0.12 ;
END V11_160x60_240V_240H

VIA V11_160x60_240V_240V
  LAYER m11 ;
    RECT -0.12 -0.054 0.12 0.054 ;
  LAYER v11 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m12 ;
    RECT -0.12 -0.068 0.12 0.068 ;
END V11_160x60_240V_240V

VIA V11_40Sx120_120H_120H
  LAYER m11 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V11_40Sx120_120H_120H

VIA V11_40Sx120_120V_120H
  LAYER m11 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V11_40Sx120_120V_120H

VIA V11_40Sx120_160H_120H
  LAYER m11 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V11_40Sx120_160H_120H

VIA V11_40Sx120_160V_120H
  LAYER m11 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V11_40Sx120_160V_120H

VIA V11_40Sx120_200H_120H
  LAYER m11 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V11_40Sx120_200H_120H

VIA V11_40Sx120_200V_120H
  LAYER m11 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V11_40Sx120_200V_120H

VIA V11_40Sx120_240H_120H
  LAYER m11 ;
    RECT -0.044 -0.12 0.044 0.12 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V11_40Sx120_240H_120H

VIA V11_40Sx120_240V_120H
  LAYER m11 ;
    RECT -0.12 -0.084 0.12 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V11_40Sx120_240V_120H

VIA V11_40Sx120_60V_120H
  LAYER m11 ;
    RECT -0.03 -0.084 0.03 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V11_40Sx120_60V_120H

VIA V11_40Sx120_90V_120H
  LAYER m11 ;
    RECT -0.045 -0.084 0.045 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V11_40Sx120_90V_120H

VIA V11_40x120_120V_120V
  LAYER m11 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V11_40x120_120V_120V

VIA V11_40x120_120V_160H
  LAYER m11 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V11_40x120_120V_160H

VIA V11_40x120_120V_160V
  LAYER m11 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V11_40x120_120V_160V

VIA V11_40x120_120V_200H
  LAYER m11 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V11_40x120_120V_200H

VIA V11_40x120_120V_200V
  LAYER m11 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V11_40x120_120V_200V

VIA V11_40x120_120V_240H
  LAYER m11 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V11_40x120_120V_240H

VIA V11_40x120_120V_240V
  LAYER m11 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.12 -0.098 0.12 0.098 ;
END V11_40x120_120V_240V

VIA V11_40x120_160H_120V
  LAYER m11 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V11_40x120_160H_120V

VIA V11_40x120_160H_160H
  LAYER m11 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V11_40x120_160H_160H

VIA V11_40x120_160H_160V
  LAYER m11 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V11_40x120_160H_160V

VIA V11_40x120_160H_200H
  LAYER m11 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V11_40x120_160H_200H

VIA V11_40x120_160H_200V
  LAYER m11 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V11_40x120_160H_200V

VIA V11_40x120_160H_240H
  LAYER m11 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V11_40x120_160H_240H

VIA V11_40x120_160H_240V
  LAYER m11 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.12 -0.098 0.12 0.098 ;
END V11_40x120_160H_240V

VIA V11_40x120_160V_120V
  LAYER m11 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V11_40x120_160V_120V

VIA V11_40x120_160V_160H
  LAYER m11 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V11_40x120_160V_160H

VIA V11_40x120_160V_160V
  LAYER m11 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V11_40x120_160V_160V

VIA V11_40x120_160V_200H
  LAYER m11 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V11_40x120_160V_200H

VIA V11_40x120_160V_200V
  LAYER m11 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V11_40x120_160V_200V

VIA V11_40x120_160V_240H
  LAYER m11 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V11_40x120_160V_240H

VIA V11_40x120_160V_240V
  LAYER m11 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.12 -0.098 0.12 0.098 ;
END V11_40x120_160V_240V

VIA V11_40x120_200H_120V
  LAYER m11 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V11_40x120_200H_120V

VIA V11_40x120_200H_160H
  LAYER m11 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V11_40x120_200H_160H

VIA V11_40x120_200H_160V
  LAYER m11 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V11_40x120_200H_160V

VIA V11_40x120_200H_200H
  LAYER m11 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V11_40x120_200H_200H

VIA V11_40x120_200H_200V
  LAYER m11 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V11_40x120_200H_200V

VIA V11_40x120_200H_240H
  LAYER m11 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V11_40x120_200H_240H

VIA V11_40x120_200H_240V
  LAYER m11 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.12 -0.098 0.12 0.098 ;
END V11_40x120_200H_240V

VIA V11_40x120_200V_120V
  LAYER m11 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V11_40x120_200V_120V

VIA V11_40x120_200V_160H
  LAYER m11 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V11_40x120_200V_160H

VIA V11_40x120_200V_160V
  LAYER m11 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V11_40x120_200V_160V

VIA V11_40x120_200V_200H
  LAYER m11 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V11_40x120_200V_200H

VIA V11_40x120_200V_200V
  LAYER m11 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V11_40x120_200V_200V

VIA V11_40x120_200V_240H
  LAYER m11 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V11_40x120_200V_240H

VIA V11_40x120_200V_240V
  LAYER m11 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.12 -0.098 0.12 0.098 ;
END V11_40x120_200V_240V

VIA V11_40x120_240H_120V
  LAYER m11 ;
    RECT -0.044 -0.12 0.044 0.12 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V11_40x120_240H_120V

VIA V11_40x120_240H_160H
  LAYER m11 ;
    RECT -0.044 -0.12 0.044 0.12 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V11_40x120_240H_160H

VIA V11_40x120_240H_160V
  LAYER m11 ;
    RECT -0.044 -0.12 0.044 0.12 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V11_40x120_240H_160V

VIA V11_40x120_240H_200H
  LAYER m11 ;
    RECT -0.044 -0.12 0.044 0.12 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V11_40x120_240H_200H

VIA V11_40x120_240H_200V
  LAYER m11 ;
    RECT -0.044 -0.12 0.044 0.12 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V11_40x120_240H_200V

VIA V11_40x120_240H_240H
  LAYER m11 ;
    RECT -0.044 -0.12 0.044 0.12 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V11_40x120_240H_240H

VIA V11_40x120_240H_240V
  LAYER m11 ;
    RECT -0.044 -0.12 0.044 0.12 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.12 -0.098 0.12 0.098 ;
END V11_40x120_240H_240V

VIA V11_40x120_240V_120V
  LAYER m11 ;
    RECT -0.12 -0.084 0.12 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V11_40x120_240V_120V

VIA V11_40x120_240V_160H
  LAYER m11 ;
    RECT -0.12 -0.084 0.12 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V11_40x120_240V_160H

VIA V11_40x120_240V_160V
  LAYER m11 ;
    RECT -0.12 -0.084 0.12 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V11_40x120_240V_160V

VIA V11_40x120_240V_200H
  LAYER m11 ;
    RECT -0.12 -0.084 0.12 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V11_40x120_240V_200H

VIA V11_40x120_240V_200V
  LAYER m11 ;
    RECT -0.12 -0.084 0.12 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V11_40x120_240V_200V

VIA V11_40x120_240V_240H
  LAYER m11 ;
    RECT -0.12 -0.084 0.12 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V11_40x120_240V_240H

VIA V11_40x120_240V_240V
  LAYER m11 ;
    RECT -0.12 -0.084 0.12 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.12 -0.098 0.12 0.098 ;
END V11_40x120_240V_240V

VIA V11_40x120_90V_120V
  LAYER m11 ;
    RECT -0.045 -0.084 0.045 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V11_40x120_90V_120V

VIA V11_40x120_90V_160H
  LAYER m11 ;
    RECT -0.045 -0.084 0.045 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V11_40x120_90V_160H

VIA V11_40x120_90V_160V
  LAYER m11 ;
    RECT -0.045 -0.084 0.045 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V11_40x120_90V_160V

VIA V11_40x120_90V_200H
  LAYER m11 ;
    RECT -0.045 -0.084 0.045 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V11_40x120_90V_200H

VIA V11_40x120_90V_200V
  LAYER m11 ;
    RECT -0.045 -0.084 0.045 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V11_40x120_90V_200V

VIA V11_40x120_90V_240H
  LAYER m11 ;
    RECT -0.045 -0.084 0.045 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.058 -0.12 0.058 0.12 ;
END V11_40x120_90V_240H

VIA V11_40x120_90V_240V
  LAYER m11 ;
    RECT -0.045 -0.084 0.045 0.084 ;
  LAYER v11 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m12 ;
    RECT -0.12 -0.098 0.12 0.098 ;
END V11_40x120_90V_240V

VIA V11_60Sx120_120H_120H
  LAYER m11 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v11 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m12 ;
    RECT -0.068 -0.06 0.068 0.06 ;
END V11_60Sx120_120H_120H

VIA V11_60Sx120_120V_120H
  LAYER m11 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v11 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m12 ;
    RECT -0.068 -0.06 0.068 0.06 ;
END V11_60Sx120_120V_120H

VIA V11_60Sx120_160H_120H
  LAYER m11 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v11 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m12 ;
    RECT -0.068 -0.06 0.068 0.06 ;
END V11_60Sx120_160H_120H

VIA V11_60Sx120_160V_120H
  LAYER m11 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v11 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m12 ;
    RECT -0.068 -0.06 0.068 0.06 ;
END V11_60Sx120_160V_120H

VIA V11_60Sx120_200H_120H
  LAYER m11 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v11 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m12 ;
    RECT -0.068 -0.06 0.068 0.06 ;
END V11_60Sx120_200H_120H

VIA V11_60Sx120_200V_120H
  LAYER m11 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v11 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m12 ;
    RECT -0.068 -0.06 0.068 0.06 ;
END V11_60Sx120_200V_120H

VIA V11_60Sx120_240H_120H
  LAYER m11 ;
    RECT -0.054 -0.12 0.054 0.12 ;
  LAYER v11 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m12 ;
    RECT -0.068 -0.06 0.068 0.06 ;
END V11_60Sx120_240H_120H

VIA V11_60Sx120_240V_120H
  LAYER m11 ;
    RECT -0.12 -0.084 0.12 0.084 ;
  LAYER v11 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m12 ;
    RECT -0.068 -0.06 0.068 0.06 ;
END V11_60Sx120_240V_120H

VIA V11_60Sx120_60V_120H
  LAYER m11 ;
    RECT -0.03 -0.084 0.03 0.084 ;
  LAYER v11 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m12 ;
    RECT -0.068 -0.06 0.068 0.06 ;
END V11_60Sx120_60V_120H

VIA V11_60Sx120_90V_120H
  LAYER m11 ;
    RECT -0.045 -0.084 0.045 0.084 ;
  LAYER v11 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m12 ;
    RECT -0.068 -0.06 0.068 0.06 ;
END V11_60Sx120_90V_120H

VIA V11_60Sx160_120V_160H
  LAYER m11 ;
    RECT -0.06 -0.104 0.06 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.08 0.068 0.08 ;
END V11_60Sx160_120V_160H

VIA V11_60Sx160_160H_160H
  LAYER m11 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.08 0.068 0.08 ;
END V11_60Sx160_160H_160H

VIA V11_60Sx160_160V_160H
  LAYER m11 ;
    RECT -0.08 -0.104 0.08 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.08 0.068 0.08 ;
END V11_60Sx160_160V_160H

VIA V11_60Sx160_200H_160H
  LAYER m11 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.08 0.068 0.08 ;
END V11_60Sx160_200H_160H

VIA V11_60Sx160_200V_160H
  LAYER m11 ;
    RECT -0.1 -0.104 0.1 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.08 0.068 0.08 ;
END V11_60Sx160_200V_160H

VIA V11_60Sx160_240H_160H
  LAYER m11 ;
    RECT -0.054 -0.12 0.054 0.12 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.08 0.068 0.08 ;
END V11_60Sx160_240H_160H

VIA V11_60Sx160_240V_160H
  LAYER m11 ;
    RECT -0.12 -0.104 0.12 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.08 0.068 0.08 ;
END V11_60Sx160_240V_160H

VIA V11_60Sx160_60V_160H
  LAYER m11 ;
    RECT -0.03 -0.104 0.03 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.08 0.068 0.08 ;
END V11_60Sx160_60V_160H

VIA V11_60Sx160_90V_160H
  LAYER m11 ;
    RECT -0.045 -0.104 0.045 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.08 0.068 0.08 ;
END V11_60Sx160_90V_160H

VIA V11_60Sx60_120H_60H
  LAYER m11 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v11 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m12 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V11_60Sx60_120H_60H

VIA V11_60Sx60_120V_60H
  LAYER m11 ;
    RECT -0.06 -0.054 0.06 0.054 ;
  LAYER v11 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m12 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V11_60Sx60_120V_60H

VIA V11_60Sx60_160H_60H
  LAYER m11 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v11 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m12 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V11_60Sx60_160H_60H

VIA V11_60Sx60_160V_60H
  LAYER m11 ;
    RECT -0.08 -0.054 0.08 0.054 ;
  LAYER v11 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m12 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V11_60Sx60_160V_60H

VIA V11_60Sx60_200H_60H
  LAYER m11 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v11 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m12 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V11_60Sx60_200H_60H

VIA V11_60Sx60_200V_60H
  LAYER m11 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v11 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m12 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V11_60Sx60_200V_60H

VIA V11_60Sx60_240H_60H
  LAYER m11 ;
    RECT -0.054 -0.12 0.054 0.12 ;
  LAYER v11 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m12 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V11_60Sx60_240H_60H

VIA V11_60Sx60_240V_60H
  LAYER m11 ;
    RECT -0.12 -0.054 0.12 0.054 ;
  LAYER v11 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m12 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V11_60Sx60_240V_60H

VIA V11_60Sx60_60V_60H
  LAYER m11 ;
    RECT -0.03 -0.054 0.03 0.054 ;
  LAYER v11 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m12 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V11_60Sx60_60V_60H

VIA V11_60Sx60_90V_60H
  LAYER m11 ;
    RECT -0.045 -0.054 0.045 0.054 ;
  LAYER v11 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m12 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V11_60Sx60_90V_60H

VIA V11_60Sx90_120H_90H
  LAYER m11 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v11 ;
    RECT -0.03 -0.045 0.03 0.045 ;
  LAYER m12 ;
    RECT -0.068 -0.045 0.068 0.045 ;
END V11_60Sx90_120H_90H

VIA V11_60Sx90_120V_90H
  LAYER m11 ;
    RECT -0.06 -0.069 0.06 0.069 ;
  LAYER v11 ;
    RECT -0.03 -0.045 0.03 0.045 ;
  LAYER m12 ;
    RECT -0.068 -0.045 0.068 0.045 ;
END V11_60Sx90_120V_90H

VIA V11_60Sx90_160H_90H
  LAYER m11 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v11 ;
    RECT -0.03 -0.045 0.03 0.045 ;
  LAYER m12 ;
    RECT -0.068 -0.045 0.068 0.045 ;
END V11_60Sx90_160H_90H

VIA V11_60Sx90_160V_90H
  LAYER m11 ;
    RECT -0.08 -0.069 0.08 0.069 ;
  LAYER v11 ;
    RECT -0.03 -0.045 0.03 0.045 ;
  LAYER m12 ;
    RECT -0.068 -0.045 0.068 0.045 ;
END V11_60Sx90_160V_90H

VIA V11_60Sx90_200H_90H
  LAYER m11 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v11 ;
    RECT -0.03 -0.045 0.03 0.045 ;
  LAYER m12 ;
    RECT -0.068 -0.045 0.068 0.045 ;
END V11_60Sx90_200H_90H

VIA V11_60Sx90_200V_90H
  LAYER m11 ;
    RECT -0.1 -0.069 0.1 0.069 ;
  LAYER v11 ;
    RECT -0.03 -0.045 0.03 0.045 ;
  LAYER m12 ;
    RECT -0.068 -0.045 0.068 0.045 ;
END V11_60Sx90_200V_90H

VIA V11_60Sx90_240H_90H
  LAYER m11 ;
    RECT -0.054 -0.12 0.054 0.12 ;
  LAYER v11 ;
    RECT -0.03 -0.045 0.03 0.045 ;
  LAYER m12 ;
    RECT -0.068 -0.045 0.068 0.045 ;
END V11_60Sx90_240H_90H

VIA V11_60Sx90_240V_90H
  LAYER m11 ;
    RECT -0.12 -0.069 0.12 0.069 ;
  LAYER v11 ;
    RECT -0.03 -0.045 0.03 0.045 ;
  LAYER m12 ;
    RECT -0.068 -0.045 0.068 0.045 ;
END V11_60Sx90_240V_90H

VIA V11_60Sx90_60V_90H
  LAYER m11 ;
    RECT -0.03 -0.069 0.03 0.069 ;
  LAYER v11 ;
    RECT -0.03 -0.045 0.03 0.045 ;
  LAYER m12 ;
    RECT -0.068 -0.045 0.068 0.045 ;
END V11_60Sx90_60V_90H

VIA V11_60Sx90_90V_90H
  LAYER m11 ;
    RECT -0.045 -0.069 0.045 0.069 ;
  LAYER v11 ;
    RECT -0.03 -0.045 0.03 0.045 ;
  LAYER m12 ;
    RECT -0.068 -0.045 0.068 0.045 ;
END V11_60Sx90_90V_90H

VIA V11_60x160_120V_120V
  LAYER m11 ;
    RECT -0.06 -0.104 0.06 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.06 -0.118 0.06 0.118 ;
END V11_60x160_120V_120V

VIA V11_60x160_120V_160V
  LAYER m11 ;
    RECT -0.06 -0.104 0.06 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.08 -0.118 0.08 0.118 ;
END V11_60x160_120V_160V

VIA V11_60x160_120V_200H
  LAYER m11 ;
    RECT -0.06 -0.104 0.06 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.1 0.068 0.1 ;
END V11_60x160_120V_200H

VIA V11_60x160_120V_200V
  LAYER m11 ;
    RECT -0.06 -0.104 0.06 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.1 -0.118 0.1 0.118 ;
END V11_60x160_120V_200V

VIA V11_60x160_120V_240H
  LAYER m11 ;
    RECT -0.06 -0.104 0.06 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.12 0.068 0.12 ;
END V11_60x160_120V_240H

VIA V11_60x160_120V_240V
  LAYER m11 ;
    RECT -0.06 -0.104 0.06 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.12 -0.118 0.12 0.118 ;
END V11_60x160_120V_240V

VIA V11_60x160_160V_120V
  LAYER m11 ;
    RECT -0.08 -0.104 0.08 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.06 -0.118 0.06 0.118 ;
END V11_60x160_160V_120V

VIA V11_60x160_160V_160V
  LAYER m11 ;
    RECT -0.08 -0.104 0.08 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.08 -0.118 0.08 0.118 ;
END V11_60x160_160V_160V

VIA V11_60x160_160V_200H
  LAYER m11 ;
    RECT -0.08 -0.104 0.08 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.1 0.068 0.1 ;
END V11_60x160_160V_200H

VIA V11_60x160_160V_200V
  LAYER m11 ;
    RECT -0.08 -0.104 0.08 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.1 -0.118 0.1 0.118 ;
END V11_60x160_160V_200V

VIA V11_60x160_160V_240H
  LAYER m11 ;
    RECT -0.08 -0.104 0.08 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.12 0.068 0.12 ;
END V11_60x160_160V_240H

VIA V11_60x160_160V_240V
  LAYER m11 ;
    RECT -0.08 -0.104 0.08 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.12 -0.118 0.12 0.118 ;
END V11_60x160_160V_240V

VIA V11_60x160_200H_120V
  LAYER m11 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.06 -0.118 0.06 0.118 ;
END V11_60x160_200H_120V

VIA V11_60x160_200H_160V
  LAYER m11 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.08 -0.118 0.08 0.118 ;
END V11_60x160_200H_160V

VIA V11_60x160_200H_200H
  LAYER m11 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.1 0.068 0.1 ;
END V11_60x160_200H_200H

VIA V11_60x160_200H_200V
  LAYER m11 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.1 -0.118 0.1 0.118 ;
END V11_60x160_200H_200V

VIA V11_60x160_200H_240H
  LAYER m11 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.12 0.068 0.12 ;
END V11_60x160_200H_240H

VIA V11_60x160_200H_240V
  LAYER m11 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.12 -0.118 0.12 0.118 ;
END V11_60x160_200H_240V

VIA V11_60x160_200V_120V
  LAYER m11 ;
    RECT -0.1 -0.104 0.1 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.06 -0.118 0.06 0.118 ;
END V11_60x160_200V_120V

VIA V11_60x160_200V_160V
  LAYER m11 ;
    RECT -0.1 -0.104 0.1 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.08 -0.118 0.08 0.118 ;
END V11_60x160_200V_160V

VIA V11_60x160_200V_200H
  LAYER m11 ;
    RECT -0.1 -0.104 0.1 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.1 0.068 0.1 ;
END V11_60x160_200V_200H

VIA V11_60x160_200V_200V
  LAYER m11 ;
    RECT -0.1 -0.104 0.1 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.1 -0.118 0.1 0.118 ;
END V11_60x160_200V_200V

VIA V11_60x160_200V_240H
  LAYER m11 ;
    RECT -0.1 -0.104 0.1 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.12 0.068 0.12 ;
END V11_60x160_200V_240H

VIA V11_60x160_200V_240V
  LAYER m11 ;
    RECT -0.1 -0.104 0.1 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.12 -0.118 0.12 0.118 ;
END V11_60x160_200V_240V

VIA V11_60x160_240H_120V
  LAYER m11 ;
    RECT -0.054 -0.12 0.054 0.12 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.06 -0.118 0.06 0.118 ;
END V11_60x160_240H_120V

VIA V11_60x160_240H_160V
  LAYER m11 ;
    RECT -0.054 -0.12 0.054 0.12 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.08 -0.118 0.08 0.118 ;
END V11_60x160_240H_160V

VIA V11_60x160_240H_200H
  LAYER m11 ;
    RECT -0.054 -0.12 0.054 0.12 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.1 0.068 0.1 ;
END V11_60x160_240H_200H

VIA V11_60x160_240H_200V
  LAYER m11 ;
    RECT -0.054 -0.12 0.054 0.12 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.1 -0.118 0.1 0.118 ;
END V11_60x160_240H_200V

VIA V11_60x160_240H_240H
  LAYER m11 ;
    RECT -0.054 -0.12 0.054 0.12 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.12 0.068 0.12 ;
END V11_60x160_240H_240H

VIA V11_60x160_240H_240V
  LAYER m11 ;
    RECT -0.054 -0.12 0.054 0.12 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.12 -0.118 0.12 0.118 ;
END V11_60x160_240H_240V

VIA V11_60x160_240V_120V
  LAYER m11 ;
    RECT -0.12 -0.104 0.12 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.06 -0.118 0.06 0.118 ;
END V11_60x160_240V_120V

VIA V11_60x160_240V_160V
  LAYER m11 ;
    RECT -0.12 -0.104 0.12 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.08 -0.118 0.08 0.118 ;
END V11_60x160_240V_160V

VIA V11_60x160_240V_200H
  LAYER m11 ;
    RECT -0.12 -0.104 0.12 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.1 0.068 0.1 ;
END V11_60x160_240V_200H

VIA V11_60x160_240V_200V
  LAYER m11 ;
    RECT -0.12 -0.104 0.12 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.1 -0.118 0.1 0.118 ;
END V11_60x160_240V_200V

VIA V11_60x160_240V_240H
  LAYER m11 ;
    RECT -0.12 -0.104 0.12 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.068 -0.12 0.068 0.12 ;
END V11_60x160_240V_240H

VIA V11_60x160_240V_240V
  LAYER m11 ;
    RECT -0.12 -0.104 0.12 0.104 ;
  LAYER v11 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m12 ;
    RECT -0.12 -0.118 0.12 0.118 ;
END V11_60x160_240V_240V

VIA V11_90Sx120_120H_120H
  LAYER m11 ;
    RECT -0.069 -0.06 0.069 0.06 ;
  LAYER v11 ;
    RECT -0.045 -0.06 0.045 0.06 ;
  LAYER m12 ;
    RECT -0.083 -0.06 0.083 0.06 ;
END V11_90Sx120_120H_120H

VIA V11_90Sx120_120V_120H
  LAYER m11 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v11 ;
    RECT -0.045 -0.06 0.045 0.06 ;
  LAYER m12 ;
    RECT -0.083 -0.06 0.083 0.06 ;
END V11_90Sx120_120V_120H

VIA V11_90Sx120_160H_120H
  LAYER m11 ;
    RECT -0.069 -0.08 0.069 0.08 ;
  LAYER v11 ;
    RECT -0.045 -0.06 0.045 0.06 ;
  LAYER m12 ;
    RECT -0.083 -0.06 0.083 0.06 ;
END V11_90Sx120_160H_120H

VIA V11_90Sx120_160V_120H
  LAYER m11 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v11 ;
    RECT -0.045 -0.06 0.045 0.06 ;
  LAYER m12 ;
    RECT -0.083 -0.06 0.083 0.06 ;
END V11_90Sx120_160V_120H

VIA V11_90Sx120_200H_120H
  LAYER m11 ;
    RECT -0.069 -0.1 0.069 0.1 ;
  LAYER v11 ;
    RECT -0.045 -0.06 0.045 0.06 ;
  LAYER m12 ;
    RECT -0.083 -0.06 0.083 0.06 ;
END V11_90Sx120_200H_120H

VIA V11_90Sx120_200V_120H
  LAYER m11 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v11 ;
    RECT -0.045 -0.06 0.045 0.06 ;
  LAYER m12 ;
    RECT -0.083 -0.06 0.083 0.06 ;
END V11_90Sx120_200V_120H

VIA V11_90Sx120_240H_120H
  LAYER m11 ;
    RECT -0.069 -0.12 0.069 0.12 ;
  LAYER v11 ;
    RECT -0.045 -0.06 0.045 0.06 ;
  LAYER m12 ;
    RECT -0.083 -0.06 0.083 0.06 ;
END V11_90Sx120_240H_120H

VIA V11_90Sx120_240V_120H
  LAYER m11 ;
    RECT -0.12 -0.084 0.12 0.084 ;
  LAYER v11 ;
    RECT -0.045 -0.06 0.045 0.06 ;
  LAYER m12 ;
    RECT -0.083 -0.06 0.083 0.06 ;
END V11_90Sx120_240V_120H

VIA V11_90Sx120_90V_120H
  LAYER m11 ;
    RECT -0.045 -0.084 0.045 0.084 ;
  LAYER v11 ;
    RECT -0.045 -0.06 0.045 0.06 ;
  LAYER m12 ;
    RECT -0.083 -0.06 0.083 0.06 ;
END V11_90Sx120_90V_120H

VIA V11_90Sx60_120H_60H
  LAYER m11 ;
    RECT -0.069 -0.06 0.069 0.06 ;
  LAYER v11 ;
    RECT -0.045 -0.03 0.045 0.03 ;
  LAYER m12 ;
    RECT -0.083 -0.03 0.083 0.03 ;
END V11_90Sx60_120H_60H

VIA V11_90Sx60_120V_60H
  LAYER m11 ;
    RECT -0.06 -0.054 0.06 0.054 ;
  LAYER v11 ;
    RECT -0.045 -0.03 0.045 0.03 ;
  LAYER m12 ;
    RECT -0.083 -0.03 0.083 0.03 ;
END V11_90Sx60_120V_60H

VIA V11_90Sx60_160H_60H
  LAYER m11 ;
    RECT -0.069 -0.08 0.069 0.08 ;
  LAYER v11 ;
    RECT -0.045 -0.03 0.045 0.03 ;
  LAYER m12 ;
    RECT -0.083 -0.03 0.083 0.03 ;
END V11_90Sx60_160H_60H

VIA V11_90Sx60_160V_60H
  LAYER m11 ;
    RECT -0.08 -0.054 0.08 0.054 ;
  LAYER v11 ;
    RECT -0.045 -0.03 0.045 0.03 ;
  LAYER m12 ;
    RECT -0.083 -0.03 0.083 0.03 ;
END V11_90Sx60_160V_60H

VIA V11_90Sx60_200H_60H
  LAYER m11 ;
    RECT -0.069 -0.1 0.069 0.1 ;
  LAYER v11 ;
    RECT -0.045 -0.03 0.045 0.03 ;
  LAYER m12 ;
    RECT -0.083 -0.03 0.083 0.03 ;
END V11_90Sx60_200H_60H

VIA V11_90Sx60_200V_60H
  LAYER m11 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v11 ;
    RECT -0.045 -0.03 0.045 0.03 ;
  LAYER m12 ;
    RECT -0.083 -0.03 0.083 0.03 ;
END V11_90Sx60_200V_60H

VIA V11_90Sx60_240H_60H
  LAYER m11 ;
    RECT -0.069 -0.12 0.069 0.12 ;
  LAYER v11 ;
    RECT -0.045 -0.03 0.045 0.03 ;
  LAYER m12 ;
    RECT -0.083 -0.03 0.083 0.03 ;
END V11_90Sx60_240H_60H

VIA V11_90Sx60_240V_60H
  LAYER m11 ;
    RECT -0.12 -0.054 0.12 0.054 ;
  LAYER v11 ;
    RECT -0.045 -0.03 0.045 0.03 ;
  LAYER m12 ;
    RECT -0.083 -0.03 0.083 0.03 ;
END V11_90Sx60_240V_60H

VIA V11_90Sx60_90V_60H
  LAYER m11 ;
    RECT -0.045 -0.054 0.045 0.054 ;
  LAYER v11 ;
    RECT -0.045 -0.03 0.045 0.03 ;
  LAYER m12 ;
    RECT -0.083 -0.03 0.083 0.03 ;
END V11_90Sx60_90V_60H

VIA V11_90Sx90_120H_90H
  LAYER m11 ;
    RECT -0.069 -0.06 0.069 0.06 ;
  LAYER v11 ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m12 ;
    RECT -0.083 -0.045 0.083 0.045 ;
END V11_90Sx90_120H_90H

VIA V11_90Sx90_120V_90H
  LAYER m11 ;
    RECT -0.06 -0.069 0.06 0.069 ;
  LAYER v11 ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m12 ;
    RECT -0.083 -0.045 0.083 0.045 ;
END V11_90Sx90_120V_90H

VIA V11_90Sx90_160H_90H
  LAYER m11 ;
    RECT -0.069 -0.08 0.069 0.08 ;
  LAYER v11 ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m12 ;
    RECT -0.083 -0.045 0.083 0.045 ;
END V11_90Sx90_160H_90H

VIA V11_90Sx90_160V_90H
  LAYER m11 ;
    RECT -0.08 -0.069 0.08 0.069 ;
  LAYER v11 ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m12 ;
    RECT -0.083 -0.045 0.083 0.045 ;
END V11_90Sx90_160V_90H

VIA V11_90Sx90_200H_90H
  LAYER m11 ;
    RECT -0.069 -0.1 0.069 0.1 ;
  LAYER v11 ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m12 ;
    RECT -0.083 -0.045 0.083 0.045 ;
END V11_90Sx90_200H_90H

VIA V11_90Sx90_200V_90H
  LAYER m11 ;
    RECT -0.1 -0.069 0.1 0.069 ;
  LAYER v11 ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m12 ;
    RECT -0.083 -0.045 0.083 0.045 ;
END V11_90Sx90_200V_90H

VIA V11_90Sx90_240H_90H
  LAYER m11 ;
    RECT -0.069 -0.12 0.069 0.12 ;
  LAYER v11 ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m12 ;
    RECT -0.083 -0.045 0.083 0.045 ;
END V11_90Sx90_240H_90H

VIA V11_90Sx90_240V_90H
  LAYER m11 ;
    RECT -0.12 -0.069 0.12 0.069 ;
  LAYER v11 ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m12 ;
    RECT -0.083 -0.045 0.083 0.045 ;
END V11_90Sx90_240V_90H

VIA V11_90Sx90_90V_90H
  LAYER m11 ;
    RECT -0.045 -0.069 0.045 0.069 ;
  LAYER v11 ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER m12 ;
    RECT -0.083 -0.045 0.083 0.045 ;
END V11_90Sx90_90V_90H

VIA V12_120x60S_120H_120V
  LAYER m12 ;
    RECT -0.104 -0.06 0.104 0.06 ;
  LAYER v12 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m13 ;
    RECT -0.06 -0.077 0.06 0.077 ;
END V12_120x60S_120H_120V

VIA V12_120x60S_120V_120V
  LAYER m12 ;
    RECT -0.06 -0.074 0.06 0.074 ;
  LAYER v12 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m13 ;
    RECT -0.06 -0.077 0.06 0.077 ;
END V12_120x60S_120V_120V

VIA V12_120x60S_160H_120V
  LAYER m12 ;
    RECT -0.104 -0.08 0.104 0.08 ;
  LAYER v12 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m13 ;
    RECT -0.06 -0.077 0.06 0.077 ;
END V12_120x60S_160H_120V

VIA V12_120x60S_160V_120V
  LAYER m12 ;
    RECT -0.08 -0.074 0.08 0.074 ;
  LAYER v12 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m13 ;
    RECT -0.06 -0.077 0.06 0.077 ;
END V12_120x60S_160V_120V

VIA V12_120x60S_200H_120V
  LAYER m12 ;
    RECT -0.104 -0.1 0.104 0.1 ;
  LAYER v12 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m13 ;
    RECT -0.06 -0.077 0.06 0.077 ;
END V12_120x60S_200H_120V

VIA V12_120x60S_200V_120V
  LAYER m12 ;
    RECT -0.1 -0.074 0.1 0.074 ;
  LAYER v12 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m13 ;
    RECT -0.06 -0.077 0.06 0.077 ;
END V12_120x60S_200V_120V

VIA V12_120x60S_240H_120V
  LAYER m12 ;
    RECT -0.104 -0.12 0.104 0.12 ;
  LAYER v12 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m13 ;
    RECT -0.06 -0.077 0.06 0.077 ;
END V12_120x60S_240H_120V

VIA V12_120x60S_240V_120V
  LAYER m12 ;
    RECT -0.12 -0.074 0.12 0.074 ;
  LAYER v12 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m13 ;
    RECT -0.06 -0.077 0.06 0.077 ;
END V12_120x60S_240V_120V

VIA V12_120x60S_60H_120V
  LAYER m12 ;
    RECT -0.104 -0.03 0.104 0.03 ;
  LAYER v12 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m13 ;
    RECT -0.06 -0.077 0.06 0.077 ;
END V12_120x60S_60H_120V

VIA V12_120x60S_90H_120V
  LAYER m12 ;
    RECT -0.104 -0.045 0.104 0.045 ;
  LAYER v12 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER m13 ;
    RECT -0.06 -0.077 0.06 0.077 ;
END V12_120x60S_90H_120V

VIA V12_160x60S_120H_160V
  LAYER m12 ;
    RECT -0.124 -0.06 0.124 0.06 ;
  LAYER v12 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m13 ;
    RECT -0.08 -0.077 0.08 0.077 ;
END V12_160x60S_120H_160V

VIA V12_160x60S_160H_160V
  LAYER m12 ;
    RECT -0.124 -0.08 0.124 0.08 ;
  LAYER v12 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m13 ;
    RECT -0.08 -0.077 0.08 0.077 ;
END V12_160x60S_160H_160V

VIA V12_160x60S_160V_160V
  LAYER m12 ;
    RECT -0.08 -0.074 0.08 0.074 ;
  LAYER v12 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m13 ;
    RECT -0.08 -0.077 0.08 0.077 ;
END V12_160x60S_160V_160V

VIA V12_160x60S_200H_160V
  LAYER m12 ;
    RECT -0.124 -0.1 0.124 0.1 ;
  LAYER v12 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m13 ;
    RECT -0.08 -0.077 0.08 0.077 ;
END V12_160x60S_200H_160V

VIA V12_160x60S_200V_160V
  LAYER m12 ;
    RECT -0.1 -0.074 0.1 0.074 ;
  LAYER v12 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m13 ;
    RECT -0.08 -0.077 0.08 0.077 ;
END V12_160x60S_200V_160V

VIA V12_160x60S_240H_160V
  LAYER m12 ;
    RECT -0.124 -0.12 0.124 0.12 ;
  LAYER v12 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m13 ;
    RECT -0.08 -0.077 0.08 0.077 ;
END V12_160x60S_240H_160V

VIA V12_160x60S_240V_160V
  LAYER m12 ;
    RECT -0.12 -0.074 0.12 0.074 ;
  LAYER v12 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m13 ;
    RECT -0.08 -0.077 0.08 0.077 ;
END V12_160x60S_240V_160V

VIA V12_160x60S_60H_160V
  LAYER m12 ;
    RECT -0.124 -0.03 0.124 0.03 ;
  LAYER v12 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m13 ;
    RECT -0.08 -0.077 0.08 0.077 ;
END V12_160x60S_60H_160V

VIA V12_160x60S_90H_160V
  LAYER m12 ;
    RECT -0.124 -0.045 0.124 0.045 ;
  LAYER v12 ;
    RECT -0.08 -0.03 0.08 0.03 ;
  LAYER m13 ;
    RECT -0.08 -0.077 0.08 0.077 ;
END V12_160x60S_90H_160V

VIA V12_240x40S_120H_240V
  LAYER m12 ;
    RECT -0.164 -0.06 0.164 0.06 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.12 -0.067 0.12 0.067 ;
END V12_240x40S_120H_240V

VIA V12_240x40S_160H_240V
  LAYER m12 ;
    RECT -0.164 -0.08 0.164 0.08 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.12 -0.067 0.12 0.067 ;
END V12_240x40S_160H_240V

VIA V12_240x40S_200H_240V
  LAYER m12 ;
    RECT -0.164 -0.1 0.164 0.1 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.12 -0.067 0.12 0.067 ;
END V12_240x40S_200H_240V

VIA V12_240x40S_240H_240V
  LAYER m12 ;
    RECT -0.164 -0.12 0.164 0.12 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.12 -0.067 0.12 0.067 ;
END V12_240x40S_240H_240V

VIA V12_240x40S_240V_240V
  LAYER m12 ;
    RECT -0.12 -0.064 0.12 0.064 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.12 -0.067 0.12 0.067 ;
END V12_240x40S_240V_240V

VIA V12_240x40S_60H_240V
  LAYER m12 ;
    RECT -0.164 -0.03 0.164 0.03 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.12 -0.067 0.12 0.067 ;
END V12_240x40S_60H_240V

VIA V12_240x40S_90H_240V
  LAYER m12 ;
    RECT -0.164 -0.045 0.164 0.045 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.12 -0.067 0.12 0.067 ;
END V12_240x40S_90H_240V

VIA V12_240x40_120H_120H
  LAYER m12 ;
    RECT -0.164 -0.06 0.164 0.06 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.06 0.167 0.06 ;
END V12_240x40_120H_120H

VIA V12_240x40_120H_160H
  LAYER m12 ;
    RECT -0.164 -0.06 0.164 0.06 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.08 0.167 0.08 ;
END V12_240x40_120H_160H

VIA V12_240x40_120H_240H
  LAYER m12 ;
    RECT -0.164 -0.06 0.164 0.06 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.12 0.167 0.12 ;
END V12_240x40_120H_240H

VIA V12_240x40_120H_320H
  LAYER m12 ;
    RECT -0.164 -0.06 0.164 0.06 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.16 0.167 0.16 ;
END V12_240x40_120H_320H

VIA V12_240x40_120H_320V
  LAYER m12 ;
    RECT -0.164 -0.06 0.164 0.06 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.16 -0.067 0.16 0.067 ;
END V12_240x40_120H_320V

VIA V12_240x40_120H_400H
  LAYER m12 ;
    RECT -0.164 -0.06 0.164 0.06 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.2 0.167 0.2 ;
END V12_240x40_120H_400H

VIA V12_240x40_120H_400V
  LAYER m12 ;
    RECT -0.164 -0.06 0.164 0.06 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.2 -0.067 0.2 0.067 ;
END V12_240x40_120H_400V

VIA V12_240x40_160H_120H
  LAYER m12 ;
    RECT -0.164 -0.08 0.164 0.08 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.06 0.167 0.06 ;
END V12_240x40_160H_120H

VIA V12_240x40_160H_160H
  LAYER m12 ;
    RECT -0.164 -0.08 0.164 0.08 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.08 0.167 0.08 ;
END V12_240x40_160H_160H

VIA V12_240x40_160H_240H
  LAYER m12 ;
    RECT -0.164 -0.08 0.164 0.08 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.12 0.167 0.12 ;
END V12_240x40_160H_240H

VIA V12_240x40_160H_320H
  LAYER m12 ;
    RECT -0.164 -0.08 0.164 0.08 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.16 0.167 0.16 ;
END V12_240x40_160H_320H

VIA V12_240x40_160H_320V
  LAYER m12 ;
    RECT -0.164 -0.08 0.164 0.08 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.16 -0.067 0.16 0.067 ;
END V12_240x40_160H_320V

VIA V12_240x40_160H_400H
  LAYER m12 ;
    RECT -0.164 -0.08 0.164 0.08 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.2 0.167 0.2 ;
END V12_240x40_160H_400H

VIA V12_240x40_160H_400V
  LAYER m12 ;
    RECT -0.164 -0.08 0.164 0.08 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.2 -0.067 0.2 0.067 ;
END V12_240x40_160H_400V

VIA V12_240x40_200H_120H
  LAYER m12 ;
    RECT -0.164 -0.1 0.164 0.1 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.06 0.167 0.06 ;
END V12_240x40_200H_120H

VIA V12_240x40_200H_160H
  LAYER m12 ;
    RECT -0.164 -0.1 0.164 0.1 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.08 0.167 0.08 ;
END V12_240x40_200H_160H

VIA V12_240x40_200H_240H
  LAYER m12 ;
    RECT -0.164 -0.1 0.164 0.1 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.12 0.167 0.12 ;
END V12_240x40_200H_240H

VIA V12_240x40_200H_320H
  LAYER m12 ;
    RECT -0.164 -0.1 0.164 0.1 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.16 0.167 0.16 ;
END V12_240x40_200H_320H

VIA V12_240x40_200H_320V
  LAYER m12 ;
    RECT -0.164 -0.1 0.164 0.1 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.16 -0.067 0.16 0.067 ;
END V12_240x40_200H_320V

VIA V12_240x40_200H_400H
  LAYER m12 ;
    RECT -0.164 -0.1 0.164 0.1 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.2 0.167 0.2 ;
END V12_240x40_200H_400H

VIA V12_240x40_200H_400V
  LAYER m12 ;
    RECT -0.164 -0.1 0.164 0.1 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.2 -0.067 0.2 0.067 ;
END V12_240x40_200H_400V

VIA V12_240x40_240H_120H
  LAYER m12 ;
    RECT -0.164 -0.12 0.164 0.12 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.06 0.167 0.06 ;
END V12_240x40_240H_120H

VIA V12_240x40_240H_160H
  LAYER m12 ;
    RECT -0.164 -0.12 0.164 0.12 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.08 0.167 0.08 ;
END V12_240x40_240H_160H

VIA V12_240x40_240H_240H
  LAYER m12 ;
    RECT -0.164 -0.12 0.164 0.12 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.12 0.167 0.12 ;
END V12_240x40_240H_240H

VIA V12_240x40_240H_320H
  LAYER m12 ;
    RECT -0.164 -0.12 0.164 0.12 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.16 0.167 0.16 ;
END V12_240x40_240H_320H

VIA V12_240x40_240H_320V
  LAYER m12 ;
    RECT -0.164 -0.12 0.164 0.12 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.16 -0.067 0.16 0.067 ;
END V12_240x40_240H_320V

VIA V12_240x40_240H_400H
  LAYER m12 ;
    RECT -0.164 -0.12 0.164 0.12 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.2 0.167 0.2 ;
END V12_240x40_240H_400H

VIA V12_240x40_240H_400V
  LAYER m12 ;
    RECT -0.164 -0.12 0.164 0.12 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.2 -0.067 0.2 0.067 ;
END V12_240x40_240H_400V

VIA V12_240x40_90H_120H
  LAYER m12 ;
    RECT -0.164 -0.045 0.164 0.045 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.06 0.167 0.06 ;
END V12_240x40_90H_120H

VIA V12_240x40_90H_160H
  LAYER m12 ;
    RECT -0.164 -0.045 0.164 0.045 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.08 0.167 0.08 ;
END V12_240x40_90H_160H

VIA V12_240x40_90H_240H
  LAYER m12 ;
    RECT -0.164 -0.045 0.164 0.045 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.12 0.167 0.12 ;
END V12_240x40_90H_240H

VIA V12_240x40_90H_320H
  LAYER m12 ;
    RECT -0.164 -0.045 0.164 0.045 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.16 0.167 0.16 ;
END V12_240x40_90H_320H

VIA V12_240x40_90H_320V
  LAYER m12 ;
    RECT -0.164 -0.045 0.164 0.045 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.16 -0.067 0.16 0.067 ;
END V12_240x40_90H_320V

VIA V12_240x40_90H_400H
  LAYER m12 ;
    RECT -0.164 -0.045 0.164 0.045 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.167 -0.2 0.167 0.2 ;
END V12_240x40_90H_400H

VIA V12_240x40_90H_400V
  LAYER m12 ;
    RECT -0.164 -0.045 0.164 0.045 ;
  LAYER v12 ;
    RECT -0.12 -0.02 0.12 0.02 ;
  LAYER m13 ;
    RECT -0.2 -0.067 0.2 0.067 ;
END V12_240x40_90H_400V

VIA V12_40Sx240_120V_240H
  LAYER m12 ;
    RECT -0.06 -0.164 0.06 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.067 -0.12 0.067 0.12 ;
END V12_40Sx240_120V_240H

VIA V12_40Sx240_160V_240H
  LAYER m12 ;
    RECT -0.08 -0.164 0.08 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.067 -0.12 0.067 0.12 ;
END V12_40Sx240_160V_240H

VIA V12_40Sx240_200V_240H
  LAYER m12 ;
    RECT -0.1 -0.164 0.1 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.067 -0.12 0.067 0.12 ;
END V12_40Sx240_200V_240H

VIA V12_40Sx240_240H_240H
  LAYER m12 ;
    RECT -0.064 -0.12 0.064 0.12 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.067 -0.12 0.067 0.12 ;
END V12_40Sx240_240H_240H

VIA V12_40Sx240_240V_240H
  LAYER m12 ;
    RECT -0.12 -0.164 0.12 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.067 -0.12 0.067 0.12 ;
END V12_40Sx240_240V_240H

VIA V12_40x240_120V_120V
  LAYER m12 ;
    RECT -0.06 -0.164 0.06 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.06 -0.167 0.06 0.167 ;
END V12_40x240_120V_120V

VIA V12_40x240_120V_160V
  LAYER m12 ;
    RECT -0.06 -0.164 0.06 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.08 -0.167 0.08 0.167 ;
END V12_40x240_120V_160V

VIA V12_40x240_120V_240V
  LAYER m12 ;
    RECT -0.06 -0.164 0.06 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.12 -0.167 0.12 0.167 ;
END V12_40x240_120V_240V

VIA V12_40x240_120V_320H
  LAYER m12 ;
    RECT -0.06 -0.164 0.06 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.067 -0.16 0.067 0.16 ;
END V12_40x240_120V_320H

VIA V12_40x240_120V_320V
  LAYER m12 ;
    RECT -0.06 -0.164 0.06 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.16 -0.167 0.16 0.167 ;
END V12_40x240_120V_320V

VIA V12_40x240_120V_400H
  LAYER m12 ;
    RECT -0.06 -0.164 0.06 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.067 -0.2 0.067 0.2 ;
END V12_40x240_120V_400H

VIA V12_40x240_120V_400V
  LAYER m12 ;
    RECT -0.06 -0.164 0.06 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.2 -0.167 0.2 0.167 ;
END V12_40x240_120V_400V

VIA V12_40x240_160V_120V
  LAYER m12 ;
    RECT -0.08 -0.164 0.08 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.06 -0.167 0.06 0.167 ;
END V12_40x240_160V_120V

VIA V12_40x240_160V_160V
  LAYER m12 ;
    RECT -0.08 -0.164 0.08 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.08 -0.167 0.08 0.167 ;
END V12_40x240_160V_160V

VIA V12_40x240_160V_240V
  LAYER m12 ;
    RECT -0.08 -0.164 0.08 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.12 -0.167 0.12 0.167 ;
END V12_40x240_160V_240V

VIA V12_40x240_160V_320H
  LAYER m12 ;
    RECT -0.08 -0.164 0.08 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.067 -0.16 0.067 0.16 ;
END V12_40x240_160V_320H

VIA V12_40x240_160V_320V
  LAYER m12 ;
    RECT -0.08 -0.164 0.08 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.16 -0.167 0.16 0.167 ;
END V12_40x240_160V_320V

VIA V12_40x240_160V_400H
  LAYER m12 ;
    RECT -0.08 -0.164 0.08 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.067 -0.2 0.067 0.2 ;
END V12_40x240_160V_400H

VIA V12_40x240_160V_400V
  LAYER m12 ;
    RECT -0.08 -0.164 0.08 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.2 -0.167 0.2 0.167 ;
END V12_40x240_160V_400V

VIA V12_40x240_200V_120V
  LAYER m12 ;
    RECT -0.1 -0.164 0.1 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.06 -0.167 0.06 0.167 ;
END V12_40x240_200V_120V

VIA V12_40x240_200V_160V
  LAYER m12 ;
    RECT -0.1 -0.164 0.1 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.08 -0.167 0.08 0.167 ;
END V12_40x240_200V_160V

VIA V12_40x240_200V_240V
  LAYER m12 ;
    RECT -0.1 -0.164 0.1 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.12 -0.167 0.12 0.167 ;
END V12_40x240_200V_240V

VIA V12_40x240_200V_320H
  LAYER m12 ;
    RECT -0.1 -0.164 0.1 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.067 -0.16 0.067 0.16 ;
END V12_40x240_200V_320H

VIA V12_40x240_200V_320V
  LAYER m12 ;
    RECT -0.1 -0.164 0.1 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.16 -0.167 0.16 0.167 ;
END V12_40x240_200V_320V

VIA V12_40x240_200V_400H
  LAYER m12 ;
    RECT -0.1 -0.164 0.1 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.067 -0.2 0.067 0.2 ;
END V12_40x240_200V_400H

VIA V12_40x240_200V_400V
  LAYER m12 ;
    RECT -0.1 -0.164 0.1 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.2 -0.167 0.2 0.167 ;
END V12_40x240_200V_400V

VIA V12_40x240_240V_120V
  LAYER m12 ;
    RECT -0.12 -0.164 0.12 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.06 -0.167 0.06 0.167 ;
END V12_40x240_240V_120V

VIA V12_40x240_240V_160V
  LAYER m12 ;
    RECT -0.12 -0.164 0.12 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.08 -0.167 0.08 0.167 ;
END V12_40x240_240V_160V

VIA V12_40x240_240V_240V
  LAYER m12 ;
    RECT -0.12 -0.164 0.12 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.12 -0.167 0.12 0.167 ;
END V12_40x240_240V_240V

VIA V12_40x240_240V_320H
  LAYER m12 ;
    RECT -0.12 -0.164 0.12 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.067 -0.16 0.067 0.16 ;
END V12_40x240_240V_320H

VIA V12_40x240_240V_320V
  LAYER m12 ;
    RECT -0.12 -0.164 0.12 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.16 -0.167 0.16 0.167 ;
END V12_40x240_240V_320V

VIA V12_40x240_240V_400H
  LAYER m12 ;
    RECT -0.12 -0.164 0.12 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.067 -0.2 0.067 0.2 ;
END V12_40x240_240V_400H

VIA V12_40x240_240V_400V
  LAYER m12 ;
    RECT -0.12 -0.164 0.12 0.164 ;
  LAYER v12 ;
    RECT -0.02 -0.12 0.02 0.12 ;
  LAYER m13 ;
    RECT -0.2 -0.167 0.2 0.167 ;
END V12_40x240_240V_400V

VIA V12_60Sx120_120H_120H
  LAYER m12 ;
    RECT -0.074 -0.06 0.074 0.06 ;
  LAYER v12 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m13 ;
    RECT -0.077 -0.06 0.077 0.06 ;
END V12_60Sx120_120H_120H

VIA V12_60Sx120_120V_120H
  LAYER m12 ;
    RECT -0.06 -0.104 0.06 0.104 ;
  LAYER v12 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m13 ;
    RECT -0.077 -0.06 0.077 0.06 ;
END V12_60Sx120_120V_120H

VIA V12_60Sx120_160H_120H
  LAYER m12 ;
    RECT -0.074 -0.08 0.074 0.08 ;
  LAYER v12 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m13 ;
    RECT -0.077 -0.06 0.077 0.06 ;
END V12_60Sx120_160H_120H

VIA V12_60Sx120_160V_120H
  LAYER m12 ;
    RECT -0.08 -0.104 0.08 0.104 ;
  LAYER v12 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m13 ;
    RECT -0.077 -0.06 0.077 0.06 ;
END V12_60Sx120_160V_120H

VIA V12_60Sx120_200H_120H
  LAYER m12 ;
    RECT -0.074 -0.1 0.074 0.1 ;
  LAYER v12 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m13 ;
    RECT -0.077 -0.06 0.077 0.06 ;
END V12_60Sx120_200H_120H

VIA V12_60Sx120_200V_120H
  LAYER m12 ;
    RECT -0.1 -0.104 0.1 0.104 ;
  LAYER v12 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m13 ;
    RECT -0.077 -0.06 0.077 0.06 ;
END V12_60Sx120_200V_120H

VIA V12_60Sx120_240H_120H
  LAYER m12 ;
    RECT -0.074 -0.12 0.074 0.12 ;
  LAYER v12 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m13 ;
    RECT -0.077 -0.06 0.077 0.06 ;
END V12_60Sx120_240H_120H

VIA V12_60Sx120_240V_120H
  LAYER m12 ;
    RECT -0.12 -0.104 0.12 0.104 ;
  LAYER v12 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER m13 ;
    RECT -0.077 -0.06 0.077 0.06 ;
END V12_60Sx120_240V_120H

VIA V12_60Sx160_120V_160H
  LAYER m12 ;
    RECT -0.06 -0.124 0.06 0.124 ;
  LAYER v12 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m13 ;
    RECT -0.077 -0.08 0.077 0.08 ;
END V12_60Sx160_120V_160H

VIA V12_60Sx160_160H_160H
  LAYER m12 ;
    RECT -0.074 -0.08 0.074 0.08 ;
  LAYER v12 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m13 ;
    RECT -0.077 -0.08 0.077 0.08 ;
END V12_60Sx160_160H_160H

VIA V12_60Sx160_160V_160H
  LAYER m12 ;
    RECT -0.08 -0.124 0.08 0.124 ;
  LAYER v12 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m13 ;
    RECT -0.077 -0.08 0.077 0.08 ;
END V12_60Sx160_160V_160H

VIA V12_60Sx160_200H_160H
  LAYER m12 ;
    RECT -0.074 -0.1 0.074 0.1 ;
  LAYER v12 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m13 ;
    RECT -0.077 -0.08 0.077 0.08 ;
END V12_60Sx160_200H_160H

VIA V12_60Sx160_200V_160H
  LAYER m12 ;
    RECT -0.1 -0.124 0.1 0.124 ;
  LAYER v12 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m13 ;
    RECT -0.077 -0.08 0.077 0.08 ;
END V12_60Sx160_200V_160H

VIA V12_60Sx160_240H_160H
  LAYER m12 ;
    RECT -0.074 -0.12 0.074 0.12 ;
  LAYER v12 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m13 ;
    RECT -0.077 -0.08 0.077 0.08 ;
END V12_60Sx160_240H_160H

VIA V12_60Sx160_240V_160H
  LAYER m12 ;
    RECT -0.12 -0.124 0.12 0.124 ;
  LAYER v12 ;
    RECT -0.03 -0.08 0.03 0.08 ;
  LAYER m13 ;
    RECT -0.077 -0.08 0.077 0.08 ;
END V12_60Sx160_240V_160H

VIA V12_60Sx80_120H_80H
  LAYER m12 ;
    RECT -0.074 -0.06 0.074 0.06 ;
  LAYER v12 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m13 ;
    RECT -0.077 -0.04 0.077 0.04 ;
END V12_60Sx80_120H_80H

VIA V12_60Sx80_120V_80H
  LAYER m12 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v12 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m13 ;
    RECT -0.077 -0.04 0.077 0.04 ;
END V12_60Sx80_120V_80H

VIA V12_60Sx80_160H_80H
  LAYER m12 ;
    RECT -0.074 -0.08 0.074 0.08 ;
  LAYER v12 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m13 ;
    RECT -0.077 -0.04 0.077 0.04 ;
END V12_60Sx80_160H_80H

VIA V12_60Sx80_160V_80H
  LAYER m12 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v12 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m13 ;
    RECT -0.077 -0.04 0.077 0.04 ;
END V12_60Sx80_160V_80H

VIA V12_60Sx80_200H_80H
  LAYER m12 ;
    RECT -0.074 -0.1 0.074 0.1 ;
  LAYER v12 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m13 ;
    RECT -0.077 -0.04 0.077 0.04 ;
END V12_60Sx80_200H_80H

VIA V12_60Sx80_200V_80H
  LAYER m12 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v12 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m13 ;
    RECT -0.077 -0.04 0.077 0.04 ;
END V12_60Sx80_200V_80H

VIA V12_60Sx80_240H_80H
  LAYER m12 ;
    RECT -0.074 -0.12 0.074 0.12 ;
  LAYER v12 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m13 ;
    RECT -0.077 -0.04 0.077 0.04 ;
END V12_60Sx80_240H_80H

VIA V12_60Sx80_240V_80H
  LAYER m12 ;
    RECT -0.12 -0.084 0.12 0.084 ;
  LAYER v12 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m13 ;
    RECT -0.077 -0.04 0.077 0.04 ;
END V12_60Sx80_240V_80H

VIA V12_60Sx80_90H_80H
  LAYER m12 ;
    RECT -0.074 -0.045 0.074 0.045 ;
  LAYER v12 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m13 ;
    RECT -0.077 -0.04 0.077 0.04 ;
END V12_60Sx80_90H_80H

VIA V12_80x60S_120H_80V
  LAYER m12 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v12 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m13 ;
    RECT -0.04 -0.077 0.04 0.077 ;
END V12_80x60S_120H_80V

VIA V12_80x60S_120V_80V
  LAYER m12 ;
    RECT -0.06 -0.074 0.06 0.074 ;
  LAYER v12 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m13 ;
    RECT -0.04 -0.077 0.04 0.077 ;
END V12_80x60S_120V_80V

VIA V12_80x60S_160H_80V
  LAYER m12 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v12 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m13 ;
    RECT -0.04 -0.077 0.04 0.077 ;
END V12_80x60S_160H_80V

VIA V12_80x60S_160V_80V
  LAYER m12 ;
    RECT -0.08 -0.074 0.08 0.074 ;
  LAYER v12 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m13 ;
    RECT -0.04 -0.077 0.04 0.077 ;
END V12_80x60S_160V_80V

VIA V12_80x60S_200H_80V
  LAYER m12 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v12 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m13 ;
    RECT -0.04 -0.077 0.04 0.077 ;
END V12_80x60S_200H_80V

VIA V12_80x60S_200V_80V
  LAYER m12 ;
    RECT -0.1 -0.074 0.1 0.074 ;
  LAYER v12 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m13 ;
    RECT -0.04 -0.077 0.04 0.077 ;
END V12_80x60S_200V_80V

VIA V12_80x60S_240H_80V
  LAYER m12 ;
    RECT -0.084 -0.12 0.084 0.12 ;
  LAYER v12 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m13 ;
    RECT -0.04 -0.077 0.04 0.077 ;
END V12_80x60S_240H_80V

VIA V12_80x60S_240V_80V
  LAYER m12 ;
    RECT -0.12 -0.074 0.12 0.074 ;
  LAYER v12 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m13 ;
    RECT -0.04 -0.077 0.04 0.077 ;
END V12_80x60S_240V_80V

VIA V12_80x60S_60H_80V
  LAYER m12 ;
    RECT -0.084 -0.03 0.084 0.03 ;
  LAYER v12 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m13 ;
    RECT -0.04 -0.077 0.04 0.077 ;
END V12_80x60S_60H_80V

VIA V12_80x60S_90H_80V
  LAYER m12 ;
    RECT -0.084 -0.045 0.084 0.045 ;
  LAYER v12 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m13 ;
    RECT -0.04 -0.077 0.04 0.077 ;
END V12_80x60S_90H_80V

VIA V12_80x90S_120H_80V
  LAYER m12 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v12 ;
    RECT -0.04 -0.045 0.04 0.045 ;
  LAYER m13 ;
    RECT -0.04 -0.092 0.04 0.092 ;
END V12_80x90S_120H_80V

VIA V12_80x90S_120V_80V
  LAYER m12 ;
    RECT -0.06 -0.089 0.06 0.089 ;
  LAYER v12 ;
    RECT -0.04 -0.045 0.04 0.045 ;
  LAYER m13 ;
    RECT -0.04 -0.092 0.04 0.092 ;
END V12_80x90S_120V_80V

VIA V12_80x90S_160H_80V
  LAYER m12 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v12 ;
    RECT -0.04 -0.045 0.04 0.045 ;
  LAYER m13 ;
    RECT -0.04 -0.092 0.04 0.092 ;
END V12_80x90S_160H_80V

VIA V12_80x90S_160V_80V
  LAYER m12 ;
    RECT -0.08 -0.089 0.08 0.089 ;
  LAYER v12 ;
    RECT -0.04 -0.045 0.04 0.045 ;
  LAYER m13 ;
    RECT -0.04 -0.092 0.04 0.092 ;
END V12_80x90S_160V_80V

VIA V12_80x90S_200H_80V
  LAYER m12 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v12 ;
    RECT -0.04 -0.045 0.04 0.045 ;
  LAYER m13 ;
    RECT -0.04 -0.092 0.04 0.092 ;
END V12_80x90S_200H_80V

VIA V12_80x90S_200V_80V
  LAYER m12 ;
    RECT -0.1 -0.089 0.1 0.089 ;
  LAYER v12 ;
    RECT -0.04 -0.045 0.04 0.045 ;
  LAYER m13 ;
    RECT -0.04 -0.092 0.04 0.092 ;
END V12_80x90S_200V_80V

VIA V12_80x90S_240H_80V
  LAYER m12 ;
    RECT -0.084 -0.12 0.084 0.12 ;
  LAYER v12 ;
    RECT -0.04 -0.045 0.04 0.045 ;
  LAYER m13 ;
    RECT -0.04 -0.092 0.04 0.092 ;
END V12_80x90S_240H_80V

VIA V12_80x90S_240V_80V
  LAYER m12 ;
    RECT -0.12 -0.089 0.12 0.089 ;
  LAYER v12 ;
    RECT -0.04 -0.045 0.04 0.045 ;
  LAYER m13 ;
    RECT -0.04 -0.092 0.04 0.092 ;
END V12_80x90S_240V_80V

VIA V12_80x90S_90H_80V
  LAYER m12 ;
    RECT -0.084 -0.045 0.084 0.045 ;
  LAYER v12 ;
    RECT -0.04 -0.045 0.04 0.045 ;
  LAYER m13 ;
    RECT -0.04 -0.092 0.04 0.092 ;
END V12_80x90S_90H_80V

VIA V13_120x80S_120H_120V
  LAYER m13 ;
    RECT -0.104 -0.06 0.104 0.06 ;
  LAYER v13 ;
    RECT -0.06 -0.04 0.06 0.04 ;
  LAYER m14 ;
    RECT -0.06 -0.087 0.06 0.087 ;
END V13_120x80S_120H_120V

VIA V13_120x80S_120V_120V
  LAYER m13 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v13 ;
    RECT -0.06 -0.04 0.06 0.04 ;
  LAYER m14 ;
    RECT -0.06 -0.087 0.06 0.087 ;
END V13_120x80S_120V_120V

VIA V13_120x80S_160H_120V
  LAYER m13 ;
    RECT -0.104 -0.08 0.104 0.08 ;
  LAYER v13 ;
    RECT -0.06 -0.04 0.06 0.04 ;
  LAYER m14 ;
    RECT -0.06 -0.087 0.06 0.087 ;
END V13_120x80S_160H_120V

VIA V13_120x80S_160V_120V
  LAYER m13 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v13 ;
    RECT -0.06 -0.04 0.06 0.04 ;
  LAYER m14 ;
    RECT -0.06 -0.087 0.06 0.087 ;
END V13_120x80S_160V_120V

VIA V13_120x80S_240H_120V
  LAYER m13 ;
    RECT -0.104 -0.12 0.104 0.12 ;
  LAYER v13 ;
    RECT -0.06 -0.04 0.06 0.04 ;
  LAYER m14 ;
    RECT -0.06 -0.087 0.06 0.087 ;
END V13_120x80S_240H_120V

VIA V13_120x80S_240V_120V
  LAYER m13 ;
    RECT -0.12 -0.084 0.12 0.084 ;
  LAYER v13 ;
    RECT -0.06 -0.04 0.06 0.04 ;
  LAYER m14 ;
    RECT -0.06 -0.087 0.06 0.087 ;
END V13_120x80S_240V_120V

VIA V13_120x80S_320H_120V
  LAYER m13 ;
    RECT -0.104 -0.16 0.104 0.16 ;
  LAYER v13 ;
    RECT -0.06 -0.04 0.06 0.04 ;
  LAYER m14 ;
    RECT -0.06 -0.087 0.06 0.087 ;
END V13_120x80S_320H_120V

VIA V13_120x80S_320V_120V
  LAYER m13 ;
    RECT -0.16 -0.084 0.16 0.084 ;
  LAYER v13 ;
    RECT -0.06 -0.04 0.06 0.04 ;
  LAYER m14 ;
    RECT -0.06 -0.087 0.06 0.087 ;
END V13_120x80S_320V_120V

VIA V13_120x80S_400H_120V
  LAYER m13 ;
    RECT -0.104 -0.2 0.104 0.2 ;
  LAYER v13 ;
    RECT -0.06 -0.04 0.06 0.04 ;
  LAYER m14 ;
    RECT -0.06 -0.087 0.06 0.087 ;
END V13_120x80S_400H_120V

VIA V13_120x80S_400V_120V
  LAYER m13 ;
    RECT -0.2 -0.084 0.2 0.084 ;
  LAYER v13 ;
    RECT -0.06 -0.04 0.06 0.04 ;
  LAYER m14 ;
    RECT -0.06 -0.087 0.06 0.087 ;
END V13_120x80S_400V_120V

VIA V13_120x80S_80H_120V
  LAYER m13 ;
    RECT -0.104 -0.04 0.104 0.04 ;
  LAYER v13 ;
    RECT -0.06 -0.04 0.06 0.04 ;
  LAYER m14 ;
    RECT -0.06 -0.087 0.06 0.087 ;
END V13_120x80S_80H_120V

VIA V13_160x80S_120H_160V
  LAYER m13 ;
    RECT -0.124 -0.06 0.124 0.06 ;
  LAYER v13 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER m14 ;
    RECT -0.08 -0.087 0.08 0.087 ;
END V13_160x80S_120H_160V

VIA V13_160x80S_160H_160V
  LAYER m13 ;
    RECT -0.124 -0.08 0.124 0.08 ;
  LAYER v13 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER m14 ;
    RECT -0.08 -0.087 0.08 0.087 ;
END V13_160x80S_160H_160V

VIA V13_160x80S_160V_160V
  LAYER m13 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v13 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER m14 ;
    RECT -0.08 -0.087 0.08 0.087 ;
END V13_160x80S_160V_160V

VIA V13_160x80S_240H_160V
  LAYER m13 ;
    RECT -0.124 -0.12 0.124 0.12 ;
  LAYER v13 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER m14 ;
    RECT -0.08 -0.087 0.08 0.087 ;
END V13_160x80S_240H_160V

VIA V13_160x80S_240V_160V
  LAYER m13 ;
    RECT -0.12 -0.084 0.12 0.084 ;
  LAYER v13 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER m14 ;
    RECT -0.08 -0.087 0.08 0.087 ;
END V13_160x80S_240V_160V

VIA V13_160x80S_320H_160V
  LAYER m13 ;
    RECT -0.124 -0.16 0.124 0.16 ;
  LAYER v13 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER m14 ;
    RECT -0.08 -0.087 0.08 0.087 ;
END V13_160x80S_320H_160V

VIA V13_160x80S_320V_160V
  LAYER m13 ;
    RECT -0.16 -0.084 0.16 0.084 ;
  LAYER v13 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER m14 ;
    RECT -0.08 -0.087 0.08 0.087 ;
END V13_160x80S_320V_160V

VIA V13_160x80S_400H_160V
  LAYER m13 ;
    RECT -0.124 -0.2 0.124 0.2 ;
  LAYER v13 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER m14 ;
    RECT -0.08 -0.087 0.08 0.087 ;
END V13_160x80S_400H_160V

VIA V13_160x80S_400V_160V
  LAYER m13 ;
    RECT -0.2 -0.084 0.2 0.084 ;
  LAYER v13 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER m14 ;
    RECT -0.08 -0.087 0.08 0.087 ;
END V13_160x80S_400V_160V

VIA V13_160x80S_80H_160V
  LAYER m13 ;
    RECT -0.124 -0.04 0.124 0.04 ;
  LAYER v13 ;
    RECT -0.08 -0.04 0.08 0.04 ;
  LAYER m14 ;
    RECT -0.08 -0.087 0.08 0.087 ;
END V13_160x80S_80H_160V

VIA V13_240x80S_120H_240V
  LAYER m13 ;
    RECT -0.164 -0.06 0.164 0.06 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.12 -0.087 0.12 0.087 ;
END V13_240x80S_120H_240V

VIA V13_240x80S_160H_240V
  LAYER m13 ;
    RECT -0.164 -0.08 0.164 0.08 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.12 -0.087 0.12 0.087 ;
END V13_240x80S_160H_240V

VIA V13_240x80S_240H_240V
  LAYER m13 ;
    RECT -0.164 -0.12 0.164 0.12 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.12 -0.087 0.12 0.087 ;
END V13_240x80S_240H_240V

VIA V13_240x80S_240V_240V
  LAYER m13 ;
    RECT -0.12 -0.084 0.12 0.084 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.12 -0.087 0.12 0.087 ;
END V13_240x80S_240V_240V

VIA V13_240x80S_320H_240V
  LAYER m13 ;
    RECT -0.164 -0.16 0.164 0.16 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.12 -0.087 0.12 0.087 ;
END V13_240x80S_320H_240V

VIA V13_240x80S_320V_240V
  LAYER m13 ;
    RECT -0.16 -0.084 0.16 0.084 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.12 -0.087 0.12 0.087 ;
END V13_240x80S_320V_240V

VIA V13_240x80S_400H_240V
  LAYER m13 ;
    RECT -0.164 -0.2 0.164 0.2 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.12 -0.087 0.12 0.087 ;
END V13_240x80S_400H_240V

VIA V13_240x80S_400V_240V
  LAYER m13 ;
    RECT -0.2 -0.084 0.2 0.084 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.12 -0.087 0.12 0.087 ;
END V13_240x80S_400V_240V

VIA V13_240x80S_80H_240V
  LAYER m13 ;
    RECT -0.164 -0.04 0.164 0.04 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.12 -0.087 0.12 0.087 ;
END V13_240x80S_80H_240V

VIA V13_240x80_160H_160H
  LAYER m13 ;
    RECT -0.164 -0.08 0.164 0.08 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.08 0.167 0.08 ;
END V13_240x80_160H_160H

VIA V13_240x80_160H_240H
  LAYER m13 ;
    RECT -0.164 -0.08 0.164 0.08 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.12 0.167 0.12 ;
END V13_240x80_160H_240H

VIA V13_240x80_160H_320H
  LAYER m13 ;
    RECT -0.164 -0.08 0.164 0.08 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.16 0.167 0.16 ;
END V13_240x80_160H_320H

VIA V13_240x80_160H_320V
  LAYER m13 ;
    RECT -0.164 -0.08 0.164 0.08 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.16 -0.087 0.16 0.087 ;
END V13_240x80_160H_320V

VIA V13_240x80_160H_400H
  LAYER m13 ;
    RECT -0.164 -0.08 0.164 0.08 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.2 0.167 0.2 ;
END V13_240x80_160H_400H

VIA V13_240x80_160H_400V
  LAYER m13 ;
    RECT -0.164 -0.08 0.164 0.08 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.2 -0.087 0.2 0.087 ;
END V13_240x80_160H_400V

VIA V13_240x80_240H_160H
  LAYER m13 ;
    RECT -0.164 -0.12 0.164 0.12 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.08 0.167 0.08 ;
END V13_240x80_240H_160H

VIA V13_240x80_240H_240H
  LAYER m13 ;
    RECT -0.164 -0.12 0.164 0.12 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.12 0.167 0.12 ;
END V13_240x80_240H_240H

VIA V13_240x80_240H_320H
  LAYER m13 ;
    RECT -0.164 -0.12 0.164 0.12 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.16 0.167 0.16 ;
END V13_240x80_240H_320H

VIA V13_240x80_240H_320V
  LAYER m13 ;
    RECT -0.164 -0.12 0.164 0.12 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.16 -0.087 0.16 0.087 ;
END V13_240x80_240H_320V

VIA V13_240x80_240H_400H
  LAYER m13 ;
    RECT -0.164 -0.12 0.164 0.12 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.2 0.167 0.2 ;
END V13_240x80_240H_400H

VIA V13_240x80_240H_400V
  LAYER m13 ;
    RECT -0.164 -0.12 0.164 0.12 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.2 -0.087 0.2 0.087 ;
END V13_240x80_240H_400V

VIA V13_240x80_320H_160H
  LAYER m13 ;
    RECT -0.164 -0.16 0.164 0.16 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.08 0.167 0.08 ;
END V13_240x80_320H_160H

VIA V13_240x80_320H_240H
  LAYER m13 ;
    RECT -0.164 -0.16 0.164 0.16 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.12 0.167 0.12 ;
END V13_240x80_320H_240H

VIA V13_240x80_320H_320H
  LAYER m13 ;
    RECT -0.164 -0.16 0.164 0.16 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.16 0.167 0.16 ;
END V13_240x80_320H_320H

VIA V13_240x80_320H_320V
  LAYER m13 ;
    RECT -0.164 -0.16 0.164 0.16 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.16 -0.087 0.16 0.087 ;
END V13_240x80_320H_320V

VIA V13_240x80_320H_400H
  LAYER m13 ;
    RECT -0.164 -0.16 0.164 0.16 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.2 0.167 0.2 ;
END V13_240x80_320H_400H

VIA V13_240x80_320H_400V
  LAYER m13 ;
    RECT -0.164 -0.16 0.164 0.16 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.2 -0.087 0.2 0.087 ;
END V13_240x80_320H_400V

VIA V13_240x80_320V_160H
  LAYER m13 ;
    RECT -0.16 -0.084 0.16 0.084 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.08 0.167 0.08 ;
END V13_240x80_320V_160H

VIA V13_240x80_320V_240H
  LAYER m13 ;
    RECT -0.16 -0.084 0.16 0.084 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.12 0.167 0.12 ;
END V13_240x80_320V_240H

VIA V13_240x80_320V_320H
  LAYER m13 ;
    RECT -0.16 -0.084 0.16 0.084 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.16 0.167 0.16 ;
END V13_240x80_320V_320H

VIA V13_240x80_320V_320V
  LAYER m13 ;
    RECT -0.16 -0.084 0.16 0.084 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.16 -0.087 0.16 0.087 ;
END V13_240x80_320V_320V

VIA V13_240x80_320V_400H
  LAYER m13 ;
    RECT -0.16 -0.084 0.16 0.084 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.2 0.167 0.2 ;
END V13_240x80_320V_400H

VIA V13_240x80_320V_400V
  LAYER m13 ;
    RECT -0.16 -0.084 0.16 0.084 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.2 -0.087 0.2 0.087 ;
END V13_240x80_320V_400V

VIA V13_240x80_400H_160H
  LAYER m13 ;
    RECT -0.164 -0.2 0.164 0.2 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.08 0.167 0.08 ;
END V13_240x80_400H_160H

VIA V13_240x80_400H_240H
  LAYER m13 ;
    RECT -0.164 -0.2 0.164 0.2 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.12 0.167 0.12 ;
END V13_240x80_400H_240H

VIA V13_240x80_400H_320H
  LAYER m13 ;
    RECT -0.164 -0.2 0.164 0.2 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.16 0.167 0.16 ;
END V13_240x80_400H_320H

VIA V13_240x80_400H_320V
  LAYER m13 ;
    RECT -0.164 -0.2 0.164 0.2 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.16 -0.087 0.16 0.087 ;
END V13_240x80_400H_320V

VIA V13_240x80_400H_400H
  LAYER m13 ;
    RECT -0.164 -0.2 0.164 0.2 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.2 0.167 0.2 ;
END V13_240x80_400H_400H

VIA V13_240x80_400H_400V
  LAYER m13 ;
    RECT -0.164 -0.2 0.164 0.2 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.2 -0.087 0.2 0.087 ;
END V13_240x80_400H_400V

VIA V13_240x80_400V_160H
  LAYER m13 ;
    RECT -0.2 -0.084 0.2 0.084 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.08 0.167 0.08 ;
END V13_240x80_400V_160H

VIA V13_240x80_400V_240H
  LAYER m13 ;
    RECT -0.2 -0.084 0.2 0.084 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.12 0.167 0.12 ;
END V13_240x80_400V_240H

VIA V13_240x80_400V_320H
  LAYER m13 ;
    RECT -0.2 -0.084 0.2 0.084 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.16 0.167 0.16 ;
END V13_240x80_400V_320H

VIA V13_240x80_400V_320V
  LAYER m13 ;
    RECT -0.2 -0.084 0.2 0.084 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.16 -0.087 0.16 0.087 ;
END V13_240x80_400V_320V

VIA V13_240x80_400V_400H
  LAYER m13 ;
    RECT -0.2 -0.084 0.2 0.084 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.167 -0.2 0.167 0.2 ;
END V13_240x80_400V_400H

VIA V13_240x80_400V_400V
  LAYER m13 ;
    RECT -0.2 -0.084 0.2 0.084 ;
  LAYER v13 ;
    RECT -0.12 -0.04 0.12 0.04 ;
  LAYER m14 ;
    RECT -0.2 -0.087 0.2 0.087 ;
END V13_240x80_400V_400V

VIA V13_80Sx120_120H_120H
  LAYER m13 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v13 ;
    RECT -0.04 -0.06 0.04 0.06 ;
  LAYER m14 ;
    RECT -0.087 -0.06 0.087 0.06 ;
END V13_80Sx120_120H_120H

VIA V13_80Sx120_120V_120H
  LAYER m13 ;
    RECT -0.06 -0.104 0.06 0.104 ;
  LAYER v13 ;
    RECT -0.04 -0.06 0.04 0.06 ;
  LAYER m14 ;
    RECT -0.087 -0.06 0.087 0.06 ;
END V13_80Sx120_120V_120H

VIA V13_80Sx120_160H_120H
  LAYER m13 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v13 ;
    RECT -0.04 -0.06 0.04 0.06 ;
  LAYER m14 ;
    RECT -0.087 -0.06 0.087 0.06 ;
END V13_80Sx120_160H_120H

VIA V13_80Sx120_160V_120H
  LAYER m13 ;
    RECT -0.08 -0.104 0.08 0.104 ;
  LAYER v13 ;
    RECT -0.04 -0.06 0.04 0.06 ;
  LAYER m14 ;
    RECT -0.087 -0.06 0.087 0.06 ;
END V13_80Sx120_160V_120H

VIA V13_80Sx120_240H_120H
  LAYER m13 ;
    RECT -0.084 -0.12 0.084 0.12 ;
  LAYER v13 ;
    RECT -0.04 -0.06 0.04 0.06 ;
  LAYER m14 ;
    RECT -0.087 -0.06 0.087 0.06 ;
END V13_80Sx120_240H_120H

VIA V13_80Sx120_240V_120H
  LAYER m13 ;
    RECT -0.12 -0.104 0.12 0.104 ;
  LAYER v13 ;
    RECT -0.04 -0.06 0.04 0.06 ;
  LAYER m14 ;
    RECT -0.087 -0.06 0.087 0.06 ;
END V13_80Sx120_240V_120H

VIA V13_80Sx120_320H_120H
  LAYER m13 ;
    RECT -0.084 -0.16 0.084 0.16 ;
  LAYER v13 ;
    RECT -0.04 -0.06 0.04 0.06 ;
  LAYER m14 ;
    RECT -0.087 -0.06 0.087 0.06 ;
END V13_80Sx120_320H_120H

VIA V13_80Sx120_320V_120H
  LAYER m13 ;
    RECT -0.16 -0.104 0.16 0.104 ;
  LAYER v13 ;
    RECT -0.04 -0.06 0.04 0.06 ;
  LAYER m14 ;
    RECT -0.087 -0.06 0.087 0.06 ;
END V13_80Sx120_320V_120H

VIA V13_80Sx120_400H_120H
  LAYER m13 ;
    RECT -0.084 -0.2 0.084 0.2 ;
  LAYER v13 ;
    RECT -0.04 -0.06 0.04 0.06 ;
  LAYER m14 ;
    RECT -0.087 -0.06 0.087 0.06 ;
END V13_80Sx120_400H_120H

VIA V13_80Sx120_400V_120H
  LAYER m13 ;
    RECT -0.2 -0.104 0.2 0.104 ;
  LAYER v13 ;
    RECT -0.04 -0.06 0.04 0.06 ;
  LAYER m14 ;
    RECT -0.087 -0.06 0.087 0.06 ;
END V13_80Sx120_400V_120H

VIA V13_80Sx120_80V_120H
  LAYER m13 ;
    RECT -0.04 -0.104 0.04 0.104 ;
  LAYER v13 ;
    RECT -0.04 -0.06 0.04 0.06 ;
  LAYER m14 ;
    RECT -0.087 -0.06 0.087 0.06 ;
END V13_80Sx120_80V_120H

VIA V13_80Sx160_120V_160H
  LAYER m13 ;
    RECT -0.06 -0.124 0.06 0.124 ;
  LAYER v13 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER m14 ;
    RECT -0.087 -0.08 0.087 0.08 ;
END V13_80Sx160_120V_160H

VIA V13_80Sx160_160H_160H
  LAYER m13 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v13 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER m14 ;
    RECT -0.087 -0.08 0.087 0.08 ;
END V13_80Sx160_160H_160H

VIA V13_80Sx160_160V_160H
  LAYER m13 ;
    RECT -0.08 -0.124 0.08 0.124 ;
  LAYER v13 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER m14 ;
    RECT -0.087 -0.08 0.087 0.08 ;
END V13_80Sx160_160V_160H

VIA V13_80Sx160_240H_160H
  LAYER m13 ;
    RECT -0.084 -0.12 0.084 0.12 ;
  LAYER v13 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER m14 ;
    RECT -0.087 -0.08 0.087 0.08 ;
END V13_80Sx160_240H_160H

VIA V13_80Sx160_240V_160H
  LAYER m13 ;
    RECT -0.12 -0.124 0.12 0.124 ;
  LAYER v13 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER m14 ;
    RECT -0.087 -0.08 0.087 0.08 ;
END V13_80Sx160_240V_160H

VIA V13_80Sx160_320H_160H
  LAYER m13 ;
    RECT -0.084 -0.16 0.084 0.16 ;
  LAYER v13 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER m14 ;
    RECT -0.087 -0.08 0.087 0.08 ;
END V13_80Sx160_320H_160H

VIA V13_80Sx160_320V_160H
  LAYER m13 ;
    RECT -0.16 -0.124 0.16 0.124 ;
  LAYER v13 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER m14 ;
    RECT -0.087 -0.08 0.087 0.08 ;
END V13_80Sx160_320V_160H

VIA V13_80Sx160_400H_160H
  LAYER m13 ;
    RECT -0.084 -0.2 0.084 0.2 ;
  LAYER v13 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER m14 ;
    RECT -0.087 -0.08 0.087 0.08 ;
END V13_80Sx160_400H_160H

VIA V13_80Sx160_400V_160H
  LAYER m13 ;
    RECT -0.2 -0.124 0.2 0.124 ;
  LAYER v13 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER m14 ;
    RECT -0.087 -0.08 0.087 0.08 ;
END V13_80Sx160_400V_160H

VIA V13_80Sx160_80V_160H
  LAYER m13 ;
    RECT -0.04 -0.124 0.04 0.124 ;
  LAYER v13 ;
    RECT -0.04 -0.08 0.04 0.08 ;
  LAYER m14 ;
    RECT -0.087 -0.08 0.087 0.08 ;
END V13_80Sx160_80V_160H

VIA V13_80Sx240_120V_240H
  LAYER m13 ;
    RECT -0.06 -0.164 0.06 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.12 0.087 0.12 ;
END V13_80Sx240_120V_240H

VIA V13_80Sx240_160V_240H
  LAYER m13 ;
    RECT -0.08 -0.164 0.08 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.12 0.087 0.12 ;
END V13_80Sx240_160V_240H

VIA V13_80Sx240_240H_240H
  LAYER m13 ;
    RECT -0.084 -0.12 0.084 0.12 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.12 0.087 0.12 ;
END V13_80Sx240_240H_240H

VIA V13_80Sx240_240V_240H
  LAYER m13 ;
    RECT -0.12 -0.164 0.12 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.12 0.087 0.12 ;
END V13_80Sx240_240V_240H

VIA V13_80Sx240_320H_240H
  LAYER m13 ;
    RECT -0.084 -0.16 0.084 0.16 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.12 0.087 0.12 ;
END V13_80Sx240_320H_240H

VIA V13_80Sx240_320V_240H
  LAYER m13 ;
    RECT -0.16 -0.164 0.16 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.12 0.087 0.12 ;
END V13_80Sx240_320V_240H

VIA V13_80Sx240_400H_240H
  LAYER m13 ;
    RECT -0.084 -0.2 0.084 0.2 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.12 0.087 0.12 ;
END V13_80Sx240_400H_240H

VIA V13_80Sx240_400V_240H
  LAYER m13 ;
    RECT -0.2 -0.164 0.2 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.12 0.087 0.12 ;
END V13_80Sx240_400V_240H

VIA V13_80Sx240_80V_240H
  LAYER m13 ;
    RECT -0.04 -0.164 0.04 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.12 0.087 0.12 ;
END V13_80Sx240_80V_240H

VIA V13_80Sx80_120H_80H
  LAYER m13 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.087 -0.04 0.087 0.04 ;
END V13_80Sx80_120H_80H

VIA V13_80Sx80_120V_80H
  LAYER m13 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.087 -0.04 0.087 0.04 ;
END V13_80Sx80_120V_80H

VIA V13_80Sx80_160H_80H
  LAYER m13 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.087 -0.04 0.087 0.04 ;
END V13_80Sx80_160H_80H

VIA V13_80Sx80_160V_80H
  LAYER m13 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.087 -0.04 0.087 0.04 ;
END V13_80Sx80_160V_80H

VIA V13_80Sx80_240H_80H
  LAYER m13 ;
    RECT -0.084 -0.12 0.084 0.12 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.087 -0.04 0.087 0.04 ;
END V13_80Sx80_240H_80H

VIA V13_80Sx80_240V_80H
  LAYER m13 ;
    RECT -0.12 -0.084 0.12 0.084 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.087 -0.04 0.087 0.04 ;
END V13_80Sx80_240V_80H

VIA V13_80Sx80_320H_80H
  LAYER m13 ;
    RECT -0.084 -0.16 0.084 0.16 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.087 -0.04 0.087 0.04 ;
END V13_80Sx80_320H_80H

VIA V13_80Sx80_320V_80H
  LAYER m13 ;
    RECT -0.16 -0.084 0.16 0.084 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.087 -0.04 0.087 0.04 ;
END V13_80Sx80_320V_80H

VIA V13_80Sx80_400H_80H
  LAYER m13 ;
    RECT -0.084 -0.2 0.084 0.2 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.087 -0.04 0.087 0.04 ;
END V13_80Sx80_400H_80H

VIA V13_80Sx80_400V_80H
  LAYER m13 ;
    RECT -0.2 -0.084 0.2 0.084 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.087 -0.04 0.087 0.04 ;
END V13_80Sx80_400V_80H

VIA V13_80Sx80_80H_80H
  LAYER m13 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.087 -0.04 0.087 0.04 ;
END V13_80Sx80_80H_80H

VIA V13_80Sx80_80V_80H
  LAYER m13 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.087 -0.04 0.087 0.04 ;
END V13_80Sx80_80V_80H

VIA V13_80x240_160V_160V
  LAYER m13 ;
    RECT -0.08 -0.164 0.08 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.08 -0.167 0.08 0.167 ;
END V13_80x240_160V_160V

VIA V13_80x240_160V_240V
  LAYER m13 ;
    RECT -0.08 -0.164 0.08 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.12 -0.167 0.12 0.167 ;
END V13_80x240_160V_240V

VIA V13_80x240_160V_320H
  LAYER m13 ;
    RECT -0.08 -0.164 0.08 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.16 0.087 0.16 ;
END V13_80x240_160V_320H

VIA V13_80x240_160V_320V
  LAYER m13 ;
    RECT -0.08 -0.164 0.08 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.16 -0.167 0.16 0.167 ;
END V13_80x240_160V_320V

VIA V13_80x240_160V_400H
  LAYER m13 ;
    RECT -0.08 -0.164 0.08 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.2 0.087 0.2 ;
END V13_80x240_160V_400H

VIA V13_80x240_160V_400V
  LAYER m13 ;
    RECT -0.08 -0.164 0.08 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.2 -0.167 0.2 0.167 ;
END V13_80x240_160V_400V

VIA V13_80x240_240V_160V
  LAYER m13 ;
    RECT -0.12 -0.164 0.12 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.08 -0.167 0.08 0.167 ;
END V13_80x240_240V_160V

VIA V13_80x240_240V_240V
  LAYER m13 ;
    RECT -0.12 -0.164 0.12 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.12 -0.167 0.12 0.167 ;
END V13_80x240_240V_240V

VIA V13_80x240_240V_320H
  LAYER m13 ;
    RECT -0.12 -0.164 0.12 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.16 0.087 0.16 ;
END V13_80x240_240V_320H

VIA V13_80x240_240V_320V
  LAYER m13 ;
    RECT -0.12 -0.164 0.12 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.16 -0.167 0.16 0.167 ;
END V13_80x240_240V_320V

VIA V13_80x240_240V_400H
  LAYER m13 ;
    RECT -0.12 -0.164 0.12 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.2 0.087 0.2 ;
END V13_80x240_240V_400H

VIA V13_80x240_240V_400V
  LAYER m13 ;
    RECT -0.12 -0.164 0.12 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.2 -0.167 0.2 0.167 ;
END V13_80x240_240V_400V

VIA V13_80x240_320H_160V
  LAYER m13 ;
    RECT -0.084 -0.16 0.084 0.16 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.08 -0.167 0.08 0.167 ;
END V13_80x240_320H_160V

VIA V13_80x240_320H_240V
  LAYER m13 ;
    RECT -0.084 -0.16 0.084 0.16 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.12 -0.167 0.12 0.167 ;
END V13_80x240_320H_240V

VIA V13_80x240_320H_320H
  LAYER m13 ;
    RECT -0.084 -0.16 0.084 0.16 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.16 0.087 0.16 ;
END V13_80x240_320H_320H

VIA V13_80x240_320H_320V
  LAYER m13 ;
    RECT -0.084 -0.16 0.084 0.16 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.16 -0.167 0.16 0.167 ;
END V13_80x240_320H_320V

VIA V13_80x240_320H_400H
  LAYER m13 ;
    RECT -0.084 -0.16 0.084 0.16 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.2 0.087 0.2 ;
END V13_80x240_320H_400H

VIA V13_80x240_320H_400V
  LAYER m13 ;
    RECT -0.084 -0.16 0.084 0.16 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.2 -0.167 0.2 0.167 ;
END V13_80x240_320H_400V

VIA V13_80x240_320V_160V
  LAYER m13 ;
    RECT -0.16 -0.164 0.16 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.08 -0.167 0.08 0.167 ;
END V13_80x240_320V_160V

VIA V13_80x240_320V_240V
  LAYER m13 ;
    RECT -0.16 -0.164 0.16 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.12 -0.167 0.12 0.167 ;
END V13_80x240_320V_240V

VIA V13_80x240_320V_320H
  LAYER m13 ;
    RECT -0.16 -0.164 0.16 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.16 0.087 0.16 ;
END V13_80x240_320V_320H

VIA V13_80x240_320V_320V
  LAYER m13 ;
    RECT -0.16 -0.164 0.16 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.16 -0.167 0.16 0.167 ;
END V13_80x240_320V_320V

VIA V13_80x240_320V_400H
  LAYER m13 ;
    RECT -0.16 -0.164 0.16 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.2 0.087 0.2 ;
END V13_80x240_320V_400H

VIA V13_80x240_320V_400V
  LAYER m13 ;
    RECT -0.16 -0.164 0.16 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.2 -0.167 0.2 0.167 ;
END V13_80x240_320V_400V

VIA V13_80x240_400H_160V
  LAYER m13 ;
    RECT -0.084 -0.2 0.084 0.2 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.08 -0.167 0.08 0.167 ;
END V13_80x240_400H_160V

VIA V13_80x240_400H_240V
  LAYER m13 ;
    RECT -0.084 -0.2 0.084 0.2 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.12 -0.167 0.12 0.167 ;
END V13_80x240_400H_240V

VIA V13_80x240_400H_320H
  LAYER m13 ;
    RECT -0.084 -0.2 0.084 0.2 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.16 0.087 0.16 ;
END V13_80x240_400H_320H

VIA V13_80x240_400H_320V
  LAYER m13 ;
    RECT -0.084 -0.2 0.084 0.2 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.16 -0.167 0.16 0.167 ;
END V13_80x240_400H_320V

VIA V13_80x240_400H_400H
  LAYER m13 ;
    RECT -0.084 -0.2 0.084 0.2 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.2 0.087 0.2 ;
END V13_80x240_400H_400H

VIA V13_80x240_400H_400V
  LAYER m13 ;
    RECT -0.084 -0.2 0.084 0.2 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.2 -0.167 0.2 0.167 ;
END V13_80x240_400H_400V

VIA V13_80x240_400V_160V
  LAYER m13 ;
    RECT -0.2 -0.164 0.2 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.08 -0.167 0.08 0.167 ;
END V13_80x240_400V_160V

VIA V13_80x240_400V_240V
  LAYER m13 ;
    RECT -0.2 -0.164 0.2 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.12 -0.167 0.12 0.167 ;
END V13_80x240_400V_240V

VIA V13_80x240_400V_320H
  LAYER m13 ;
    RECT -0.2 -0.164 0.2 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.16 0.087 0.16 ;
END V13_80x240_400V_320H

VIA V13_80x240_400V_320V
  LAYER m13 ;
    RECT -0.2 -0.164 0.2 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.16 -0.167 0.16 0.167 ;
END V13_80x240_400V_320V

VIA V13_80x240_400V_400H
  LAYER m13 ;
    RECT -0.2 -0.164 0.2 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.087 -0.2 0.087 0.2 ;
END V13_80x240_400V_400H

VIA V13_80x240_400V_400V
  LAYER m13 ;
    RECT -0.2 -0.164 0.2 0.164 ;
  LAYER v13 ;
    RECT -0.04 -0.12 0.04 0.12 ;
  LAYER m14 ;
    RECT -0.2 -0.167 0.2 0.167 ;
END V13_80x240_400V_400V

VIA V13_80x80S_120H_80V
  LAYER m13 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.04 -0.087 0.04 0.087 ;
END V13_80x80S_120H_80V

VIA V13_80x80S_120V_80V
  LAYER m13 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.04 -0.087 0.04 0.087 ;
END V13_80x80S_120V_80V

VIA V13_80x80S_160H_80V
  LAYER m13 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.04 -0.087 0.04 0.087 ;
END V13_80x80S_160H_80V

VIA V13_80x80S_160V_80V
  LAYER m13 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.04 -0.087 0.04 0.087 ;
END V13_80x80S_160V_80V

VIA V13_80x80S_240H_80V
  LAYER m13 ;
    RECT -0.084 -0.12 0.084 0.12 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.04 -0.087 0.04 0.087 ;
END V13_80x80S_240H_80V

VIA V13_80x80S_240V_80V
  LAYER m13 ;
    RECT -0.12 -0.084 0.12 0.084 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.04 -0.087 0.04 0.087 ;
END V13_80x80S_240V_80V

VIA V13_80x80S_320H_80V
  LAYER m13 ;
    RECT -0.084 -0.16 0.084 0.16 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.04 -0.087 0.04 0.087 ;
END V13_80x80S_320H_80V

VIA V13_80x80S_320V_80V
  LAYER m13 ;
    RECT -0.16 -0.084 0.16 0.084 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.04 -0.087 0.04 0.087 ;
END V13_80x80S_320V_80V

VIA V13_80x80S_400H_80V
  LAYER m13 ;
    RECT -0.084 -0.2 0.084 0.2 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.04 -0.087 0.04 0.087 ;
END V13_80x80S_400H_80V

VIA V13_80x80S_400V_80V
  LAYER m13 ;
    RECT -0.2 -0.084 0.2 0.084 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.04 -0.087 0.04 0.087 ;
END V13_80x80S_400V_80V

VIA V13_80x80S_80H_80V
  LAYER m13 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.04 -0.087 0.04 0.087 ;
END V13_80x80S_80H_80V

VIA V13_80x80S_80V_80V
  LAYER m13 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v13 ;
    RECT -0.04 -0.04 0.04 0.04 ;
  LAYER m14 ;
    RECT -0.04 -0.087 0.04 0.087 ;
END V13_80x80S_80V_80V

VIA V1_30x20_30V_20H
  LAYER m1 ;
    RECT -0.015 -0.021 0.015 0.021 ;
  LAYER v1 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m2 ;
    RECT -0.0325 -0.01 0.0325 0.01 ;
END V1_30x20_30V_20H

VIA V1_30x20_35H_20H
  LAYER m1 ;
    RECT -0.03 -0.0175 0.03 0.0175 ;
  LAYER v1 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m2 ;
    RECT -0.0325 -0.01 0.0325 0.01 ;
END V1_30x20_35H_20H

VIA V1_30x20_56H_20H
  LAYER m1 ;
    RECT -0.03 -0.028 0.03 0.028 ;
  LAYER v1 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m2 ;
    RECT -0.0325 -0.01 0.0325 0.01 ;
END V1_30x20_56H_20H

VIA V1_30x20_56V_20H
  LAYER m1 ;
    RECT -0.028 -0.021 0.028 0.021 ;
  LAYER v1 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m2 ;
    RECT -0.0325 -0.01 0.0325 0.01 ;
END V1_30x20_56V_20H

VIA V1_30x20_70V_20H
  LAYER m1 ;
    RECT -0.035 -0.021 0.035 0.021 ;
  LAYER v1 ;
    RECT -0.015 -0.01 0.015 0.01 ;
  LAYER m2 ;
    RECT -0.0325 -0.01 0.0325 0.01 ;
END V1_30x20_70V_20H

VIA V1_30x28_30V_28H
  LAYER m1 ;
    RECT -0.015 -0.025 0.015 0.025 ;
  LAYER v1 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m2 ;
    RECT -0.0325 -0.014 0.0325 0.014 ;
END V1_30x28_30V_28H

VIA V1_30x28_56H_28H
  LAYER m1 ;
    RECT -0.03 -0.028 0.03 0.028 ;
  LAYER v1 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m2 ;
    RECT -0.0325 -0.014 0.0325 0.014 ;
END V1_30x28_56H_28H

VIA V1_30x28_56V_28H
  LAYER m1 ;
    RECT -0.028 -0.025 0.028 0.025 ;
  LAYER v1 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m2 ;
    RECT -0.0325 -0.014 0.0325 0.014 ;
END V1_30x28_56V_28H

VIA V1_30x28_70V_28H
  LAYER m1 ;
    RECT -0.035 -0.025 0.035 0.025 ;
  LAYER v1 ;
    RECT -0.015 -0.014 0.015 0.014 ;
  LAYER m2 ;
    RECT -0.0325 -0.014 0.0325 0.014 ;
END V1_30x28_70V_28H

VIA V1_30x38_30V_38H
  LAYER m1 ;
    RECT -0.015 -0.03 0.015 0.03 ;
  LAYER v1 ;
    RECT -0.015 -0.019 0.015 0.019 ;
  LAYER m2 ;
    RECT -0.0325 -0.019 0.0325 0.019 ;
END V1_30x38_30V_38H

VIA V1_30x38_56H_38H
  LAYER m1 ;
    RECT -0.03 -0.028 0.03 0.028 ;
  LAYER v1 ;
    RECT -0.015 -0.019 0.015 0.019 ;
  LAYER m2 ;
    RECT -0.0325 -0.019 0.0325 0.019 ;
END V1_30x38_56H_38H

VIA V1_30x38_56V_38H
  LAYER m1 ;
    RECT -0.028 -0.03 0.028 0.03 ;
  LAYER v1 ;
    RECT -0.015 -0.019 0.015 0.019 ;
  LAYER m2 ;
    RECT -0.0325 -0.019 0.0325 0.019 ;
END V1_30x38_56V_38H

VIA V1_30x38_70V_38H
  LAYER m1 ;
    RECT -0.035 -0.03 0.035 0.03 ;
  LAYER v1 ;
    RECT -0.015 -0.019 0.015 0.019 ;
  LAYER m2 ;
    RECT -0.0325 -0.019 0.0325 0.019 ;
END V1_30x38_70V_38H

VIA V1_30x56_30V_56H
  LAYER m1 ;
    RECT -0.015 -0.039 0.015 0.039 ;
  LAYER v1 ;
    RECT -0.015 -0.028 0.015 0.028 ;
  LAYER m2 ;
    RECT -0.0325 -0.028 0.0325 0.028 ;
END V1_30x56_30V_56H

VIA V1_30x56_56H_56H
  LAYER m1 ;
    RECT -0.03 -0.028 0.03 0.028 ;
  LAYER v1 ;
    RECT -0.015 -0.028 0.015 0.028 ;
  LAYER m2 ;
    RECT -0.0325 -0.028 0.0325 0.028 ;
END V1_30x56_56H_56H

VIA V1_30x56_56V_56H
  LAYER m1 ;
    RECT -0.028 -0.039 0.028 0.039 ;
  LAYER v1 ;
    RECT -0.015 -0.028 0.015 0.028 ;
  LAYER m2 ;
    RECT -0.0325 -0.028 0.0325 0.028 ;
END V1_30x56_56V_56H

VIA V1_30x56_70V_56H
  LAYER m1 ;
    RECT -0.035 -0.039 0.035 0.039 ;
  LAYER v1 ;
    RECT -0.015 -0.028 0.015 0.028 ;
  LAYER m2 ;
    RECT -0.0325 -0.028 0.0325 0.028 ;
END V1_30x56_70V_56H

VIA V1_35x35_35H_56H
  LAYER m1 ;
    RECT -0.0325 -0.0175 0.0325 0.0175 ;
  LAYER v1 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m2 ;
    RECT -0.0225 -0.028 0.0225 0.028 ;
END V1_35x35_35H_56H

VIA V1_35x35_35H_56V
  LAYER m1 ;
    RECT -0.0325 -0.0175 0.0325 0.0175 ;
  LAYER v1 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m2 ;
    RECT -0.028 -0.0225 0.028 0.0225 ;
END V1_35x35_35H_56V

VIA V1_35x35_56H_56H
  LAYER m1 ;
    RECT -0.0325 -0.028 0.0325 0.028 ;
  LAYER v1 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m2 ;
    RECT -0.0225 -0.028 0.0225 0.028 ;
END V1_35x35_56H_56H

VIA V1_35x35_56H_56V
  LAYER m1 ;
    RECT -0.0325 -0.028 0.0325 0.028 ;
  LAYER v1 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m2 ;
    RECT -0.028 -0.0225 0.028 0.0225 ;
END V1_35x35_56H_56V

VIA V1_35x35_56V_56H
  LAYER m1 ;
    RECT -0.028 -0.0285 0.028 0.0285 ;
  LAYER v1 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m2 ;
    RECT -0.0225 -0.028 0.0225 0.028 ;
END V1_35x35_56V_56H

VIA V1_35x35_56V_56V
  LAYER m1 ;
    RECT -0.028 -0.0285 0.028 0.0285 ;
  LAYER v1 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m2 ;
    RECT -0.028 -0.0225 0.028 0.0225 ;
END V1_35x35_56V_56V

VIA V1_35x35_70V_56H
  LAYER m1 ;
    RECT -0.035 -0.0285 0.035 0.0285 ;
  LAYER v1 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m2 ;
    RECT -0.0225 -0.028 0.0225 0.028 ;
END V1_35x35_70V_56H

VIA V1_35x35_70V_56V
  LAYER m1 ;
    RECT -0.035 -0.0285 0.035 0.0285 ;
  LAYER v1 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m2 ;
    RECT -0.028 -0.0225 0.028 0.0225 ;
END V1_35x35_70V_56V

VIA V2_24x20_20H_24V
  LAYER m2 ;
    RECT -0.032 -0.01 0.032 0.01 ;
  LAYER v2 ;
    RECT -0.012 -0.01 0.012 0.01 ;
  LAYER m3 ;
    RECT -0.012 -0.034 0.012 0.034 ;
END V2_24x20_20H_24V

VIA V2_24x20_28H_24V
  LAYER m2 ;
    RECT -0.032 -0.014 0.032 0.014 ;
  LAYER v2 ;
    RECT -0.012 -0.01 0.012 0.01 ;
  LAYER m3 ;
    RECT -0.012 -0.034 0.012 0.034 ;
END V2_24x20_28H_24V

VIA V2_24x20_38H_24V
  LAYER m2 ;
    RECT -0.032 -0.019 0.032 0.019 ;
  LAYER v2 ;
    RECT -0.012 -0.01 0.012 0.01 ;
  LAYER m3 ;
    RECT -0.012 -0.034 0.012 0.034 ;
END V2_24x20_38H_24V

VIA V2_24x20_56H_24V
  LAYER m2 ;
    RECT -0.032 -0.028 0.032 0.028 ;
  LAYER v2 ;
    RECT -0.012 -0.01 0.012 0.01 ;
  LAYER m3 ;
    RECT -0.012 -0.034 0.012 0.034 ;
END V2_24x20_56H_24V

VIA V2_24x20_56V_24V
  LAYER m2 ;
    RECT -0.028 -0.03 0.028 0.03 ;
  LAYER v2 ;
    RECT -0.012 -0.01 0.012 0.01 ;
  LAYER m3 ;
    RECT -0.012 -0.034 0.012 0.034 ;
END V2_24x20_56V_24V

VIA V2_34x20_20H_34V
  LAYER m2 ;
    RECT -0.037 -0.01 0.037 0.01 ;
  LAYER v2 ;
    RECT -0.017 -0.01 0.017 0.01 ;
  LAYER m3 ;
    RECT -0.017 -0.034 0.017 0.034 ;
END V2_34x20_20H_34V

VIA V2_34x20_28H_34V
  LAYER m2 ;
    RECT -0.037 -0.014 0.037 0.014 ;
  LAYER v2 ;
    RECT -0.017 -0.01 0.017 0.01 ;
  LAYER m3 ;
    RECT -0.017 -0.034 0.017 0.034 ;
END V2_34x20_28H_34V

VIA V2_34x20_38H_34V
  LAYER m2 ;
    RECT -0.037 -0.019 0.037 0.019 ;
  LAYER v2 ;
    RECT -0.017 -0.01 0.017 0.01 ;
  LAYER m3 ;
    RECT -0.017 -0.034 0.017 0.034 ;
END V2_34x20_38H_34V

VIA V2_34x20_56H_34V
  LAYER m2 ;
    RECT -0.037 -0.028 0.037 0.028 ;
  LAYER v2 ;
    RECT -0.017 -0.01 0.017 0.01 ;
  LAYER m3 ;
    RECT -0.017 -0.034 0.017 0.034 ;
END V2_34x20_56H_34V

VIA V2_34x20_56V_34V
  LAYER m2 ;
    RECT -0.028 -0.03 0.028 0.03 ;
  LAYER v2 ;
    RECT -0.017 -0.01 0.017 0.01 ;
  LAYER m3 ;
    RECT -0.017 -0.034 0.017 0.034 ;
END V2_34x20_56V_34V

VIA V2_34x28_28H_34V
  LAYER m2 ;
    RECT -0.037 -0.014 0.037 0.014 ;
  LAYER v2 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER m3 ;
    RECT -0.017 -0.038 0.017 0.038 ;
END V2_34x28_28H_34V

VIA V2_34x28_38H_34V
  LAYER m2 ;
    RECT -0.037 -0.019 0.037 0.019 ;
  LAYER v2 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER m3 ;
    RECT -0.017 -0.038 0.017 0.038 ;
END V2_34x28_38H_34V

VIA V2_34x28_56H_34V
  LAYER m2 ;
    RECT -0.037 -0.028 0.037 0.028 ;
  LAYER v2 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER m3 ;
    RECT -0.017 -0.038 0.017 0.038 ;
END V2_34x28_56H_34V

VIA V2_34x28_56V_34V
  LAYER m2 ;
    RECT -0.028 -0.034 0.028 0.034 ;
  LAYER v2 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER m3 ;
    RECT -0.017 -0.038 0.017 0.038 ;
END V2_34x28_56V_34V

VIA V2_35x35_38H_44V
  LAYER m2 ;
    RECT -0.0375 -0.019 0.0375 0.019 ;
  LAYER v2 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m3 ;
    RECT -0.022 -0.0415 0.022 0.0415 ;
END V2_35x35_38H_44V

VIA V2_35x35_38H_56H
  LAYER m2 ;
    RECT -0.0375 -0.019 0.0375 0.019 ;
  LAYER v2 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m3 ;
    RECT -0.0415 -0.028 0.0415 0.028 ;
END V2_35x35_38H_56H

VIA V2_35x35_38H_56V
  LAYER m2 ;
    RECT -0.0375 -0.019 0.0375 0.019 ;
  LAYER v2 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m3 ;
    RECT -0.028 -0.0415 0.028 0.0415 ;
END V2_35x35_38H_56V

VIA V2_35x35_56H_44V
  LAYER m2 ;
    RECT -0.0375 -0.028 0.0375 0.028 ;
  LAYER v2 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m3 ;
    RECT -0.022 -0.0415 0.022 0.0415 ;
END V2_35x35_56H_44V

VIA V2_35x35_56H_56H
  LAYER m2 ;
    RECT -0.0375 -0.028 0.0375 0.028 ;
  LAYER v2 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m3 ;
    RECT -0.0415 -0.028 0.0415 0.028 ;
END V2_35x35_56H_56H

VIA V2_35x35_56H_56V
  LAYER m2 ;
    RECT -0.0375 -0.028 0.0375 0.028 ;
  LAYER v2 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m3 ;
    RECT -0.028 -0.0415 0.028 0.0415 ;
END V2_35x35_56H_56V

VIA V2_35x35_56V_44V
  LAYER m2 ;
    RECT -0.028 -0.0375 0.028 0.0375 ;
  LAYER v2 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m3 ;
    RECT -0.022 -0.0415 0.022 0.0415 ;
END V2_35x35_56V_44V

VIA V2_35x35_56V_56H
  LAYER m2 ;
    RECT -0.028 -0.0375 0.028 0.0375 ;
  LAYER v2 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m3 ;
    RECT -0.0415 -0.028 0.0415 0.028 ;
END V2_35x35_56V_56H

VIA V2_35x35_56V_56V
  LAYER m2 ;
    RECT -0.028 -0.0375 0.028 0.0375 ;
  LAYER v2 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m3 ;
    RECT -0.028 -0.0415 0.028 0.0415 ;
END V2_35x35_56V_56V

VIA V2_44x20_20H_44V
  LAYER m2 ;
    RECT -0.0325 -0.01 0.0325 0.01 ;
  LAYER v2 ;
    RECT -0.022 -0.01 0.022 0.01 ;
  LAYER m3 ;
    RECT -0.022 -0.034 0.022 0.034 ;
END V2_44x20_20H_44V

VIA V2_44x20_28H_44V
  LAYER m2 ;
    RECT -0.0325 -0.014 0.0325 0.014 ;
  LAYER v2 ;
    RECT -0.022 -0.01 0.022 0.01 ;
  LAYER m3 ;
    RECT -0.022 -0.034 0.022 0.034 ;
END V2_44x20_28H_44V

VIA V2_44x20_38H_44V
  LAYER m2 ;
    RECT -0.0325 -0.019 0.0325 0.019 ;
  LAYER v2 ;
    RECT -0.022 -0.01 0.022 0.01 ;
  LAYER m3 ;
    RECT -0.022 -0.034 0.022 0.034 ;
END V2_44x20_38H_44V

VIA V2_44x20_56H_44V
  LAYER m2 ;
    RECT -0.0325 -0.028 0.0325 0.028 ;
  LAYER v2 ;
    RECT -0.022 -0.01 0.022 0.01 ;
  LAYER m3 ;
    RECT -0.022 -0.034 0.022 0.034 ;
END V2_44x20_56H_44V

VIA V2_44x20_56V_44V
  LAYER m2 ;
    RECT -0.028 -0.03 0.028 0.03 ;
  LAYER v2 ;
    RECT -0.022 -0.01 0.022 0.01 ;
  LAYER m3 ;
    RECT -0.022 -0.034 0.022 0.034 ;
END V2_44x20_56V_44V

VIA V2_44x38_38H_44V
  LAYER m2 ;
    RECT -0.042 -0.019 0.042 0.019 ;
  LAYER v2 ;
    RECT -0.022 -0.019 0.022 0.019 ;
  LAYER m3 ;
    RECT -0.022 -0.043 0.022 0.043 ;
END V2_44x38_38H_44V

VIA V2_44x38_56H_44V
  LAYER m2 ;
    RECT -0.042 -0.028 0.042 0.028 ;
  LAYER v2 ;
    RECT -0.022 -0.019 0.022 0.019 ;
  LAYER m3 ;
    RECT -0.022 -0.043 0.022 0.043 ;
END V2_44x38_56H_44V

VIA V2_44x38_56V_44V
  LAYER m2 ;
    RECT -0.028 -0.039 0.028 0.039 ;
  LAYER v2 ;
    RECT -0.022 -0.019 0.022 0.019 ;
  LAYER m3 ;
    RECT -0.022 -0.043 0.022 0.043 ;
END V2_44x38_56V_44V

VIA V2_56x20_20H_56V
  LAYER m2 ;
    RECT -0.048 -0.01 0.048 0.01 ;
  LAYER v2 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m3 ;
    RECT -0.028 -0.034 0.028 0.034 ;
END V2_56x20_20H_56V

VIA V2_56x20_28H_56V
  LAYER m2 ;
    RECT -0.048 -0.014 0.048 0.014 ;
  LAYER v2 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m3 ;
    RECT -0.028 -0.034 0.028 0.034 ;
END V2_56x20_28H_56V

VIA V2_56x20_38H_56V
  LAYER m2 ;
    RECT -0.048 -0.019 0.048 0.019 ;
  LAYER v2 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m3 ;
    RECT -0.028 -0.034 0.028 0.034 ;
END V2_56x20_38H_56V

VIA V2_56x20_56H_56V
  LAYER m2 ;
    RECT -0.048 -0.028 0.048 0.028 ;
  LAYER v2 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m3 ;
    RECT -0.028 -0.034 0.028 0.034 ;
END V2_56x20_56H_56V

VIA V2_56x20_56V_56V
  LAYER m2 ;
    RECT -0.028 -0.03 0.028 0.03 ;
  LAYER v2 ;
    RECT -0.028 -0.01 0.028 0.01 ;
  LAYER m3 ;
    RECT -0.028 -0.034 0.028 0.034 ;
END V2_56x20_56V_56V

VIA V3_24x24_24V_24H
  LAYER m3 ;
    RECT -0.012 -0.036 0.012 0.036 ;
  LAYER v3 ;
    RECT -0.012 -0.012 0.012 0.012 ;
  LAYER m4 ;
    RECT -0.036 -0.012 0.036 0.012 ;
END V3_24x24_24V_24H

VIA V3_24x24_34V_24H
  LAYER m3 ;
    RECT -0.017 -0.036 0.017 0.036 ;
  LAYER v3 ;
    RECT -0.012 -0.012 0.012 0.012 ;
  LAYER m4 ;
    RECT -0.036 -0.012 0.036 0.012 ;
END V3_24x24_34V_24H

VIA V3_24x24_44V_24H
  LAYER m3 ;
    RECT -0.022 -0.036 0.022 0.036 ;
  LAYER v3 ;
    RECT -0.012 -0.012 0.012 0.012 ;
  LAYER m4 ;
    RECT -0.036 -0.012 0.036 0.012 ;
END V3_24x24_44V_24H

VIA V3_24x24_56H_24H
  LAYER m3 ;
    RECT -0.036 -0.028 0.036 0.028 ;
  LAYER v3 ;
    RECT -0.012 -0.012 0.012 0.012 ;
  LAYER m4 ;
    RECT -0.036 -0.012 0.036 0.012 ;
END V3_24x24_56H_24H

VIA V3_24x24_56V_24H
  LAYER m3 ;
    RECT -0.028 -0.036 0.028 0.036 ;
  LAYER v3 ;
    RECT -0.012 -0.012 0.012 0.012 ;
  LAYER m4 ;
    RECT -0.036 -0.012 0.036 0.012 ;
END V3_24x24_56V_24H

VIA V3_24x28_24V_28H
  LAYER m3 ;
    RECT -0.012 -0.038 0.012 0.038 ;
  LAYER v3 ;
    RECT -0.012 -0.014 0.012 0.014 ;
  LAYER m4 ;
    RECT -0.036 -0.014 0.036 0.014 ;
END V3_24x28_24V_28H

VIA V3_24x28_34V_28H
  LAYER m3 ;
    RECT -0.017 -0.038 0.017 0.038 ;
  LAYER v3 ;
    RECT -0.012 -0.014 0.012 0.014 ;
  LAYER m4 ;
    RECT -0.036 -0.014 0.036 0.014 ;
END V3_24x28_34V_28H

VIA V3_24x28_44V_28H
  LAYER m3 ;
    RECT -0.022 -0.038 0.022 0.038 ;
  LAYER v3 ;
    RECT -0.012 -0.014 0.012 0.014 ;
  LAYER m4 ;
    RECT -0.036 -0.014 0.036 0.014 ;
END V3_24x28_44V_28H

VIA V3_24x28_56H_28H
  LAYER m3 ;
    RECT -0.036 -0.028 0.036 0.028 ;
  LAYER v3 ;
    RECT -0.012 -0.014 0.012 0.014 ;
  LAYER m4 ;
    RECT -0.036 -0.014 0.036 0.014 ;
END V3_24x28_56H_28H

VIA V3_24x28_56V_28H
  LAYER m3 ;
    RECT -0.028 -0.038 0.028 0.038 ;
  LAYER v3 ;
    RECT -0.012 -0.014 0.012 0.014 ;
  LAYER m4 ;
    RECT -0.036 -0.014 0.036 0.014 ;
END V3_24x28_56V_28H

VIA V3_24x44_24V_44H
  LAYER m3 ;
    RECT -0.012 -0.046 0.012 0.046 ;
  LAYER v3 ;
    RECT -0.012 -0.022 0.012 0.022 ;
  LAYER m4 ;
    RECT -0.036 -0.022 0.036 0.022 ;
END V3_24x44_24V_44H

VIA V3_24x44_34V_44H
  LAYER m3 ;
    RECT -0.017 -0.046 0.017 0.046 ;
  LAYER v3 ;
    RECT -0.012 -0.022 0.012 0.022 ;
  LAYER m4 ;
    RECT -0.036 -0.022 0.036 0.022 ;
END V3_24x44_34V_44H

VIA V3_24x44_44V_44H
  LAYER m3 ;
    RECT -0.022 -0.046 0.022 0.046 ;
  LAYER v3 ;
    RECT -0.012 -0.022 0.012 0.022 ;
  LAYER m4 ;
    RECT -0.036 -0.022 0.036 0.022 ;
END V3_24x44_44V_44H

VIA V3_24x44_56H_44H
  LAYER m3 ;
    RECT -0.036 -0.028 0.036 0.028 ;
  LAYER v3 ;
    RECT -0.012 -0.022 0.012 0.022 ;
  LAYER m4 ;
    RECT -0.036 -0.022 0.036 0.022 ;
END V3_24x44_56H_44H

VIA V3_24x44_56V_44H
  LAYER m3 ;
    RECT -0.028 -0.046 0.028 0.046 ;
  LAYER v3 ;
    RECT -0.012 -0.022 0.012 0.022 ;
  LAYER m4 ;
    RECT -0.036 -0.022 0.036 0.022 ;
END V3_24x44_56V_44H

VIA V3_24x56_24V_56H
  LAYER m3 ;
    RECT -0.012 -0.052 0.012 0.052 ;
  LAYER v3 ;
    RECT -0.012 -0.028 0.012 0.028 ;
  LAYER m4 ;
    RECT -0.036 -0.028 0.036 0.028 ;
END V3_24x56_24V_56H

VIA V3_24x56_34V_56H
  LAYER m3 ;
    RECT -0.017 -0.052 0.017 0.052 ;
  LAYER v3 ;
    RECT -0.012 -0.028 0.012 0.028 ;
  LAYER m4 ;
    RECT -0.036 -0.028 0.036 0.028 ;
END V3_24x56_34V_56H

VIA V3_24x56_44V_56H
  LAYER m3 ;
    RECT -0.022 -0.052 0.022 0.052 ;
  LAYER v3 ;
    RECT -0.012 -0.028 0.012 0.028 ;
  LAYER m4 ;
    RECT -0.036 -0.028 0.036 0.028 ;
END V3_24x56_44V_56H

VIA V3_24x56_56H_56H
  LAYER m3 ;
    RECT -0.036 -0.028 0.036 0.028 ;
  LAYER v3 ;
    RECT -0.012 -0.028 0.012 0.028 ;
  LAYER m4 ;
    RECT -0.036 -0.028 0.036 0.028 ;
END V3_24x56_56H_56H

VIA V3_24x56_56V_56H
  LAYER m3 ;
    RECT -0.028 -0.052 0.028 0.052 ;
  LAYER v3 ;
    RECT -0.012 -0.028 0.012 0.028 ;
  LAYER m4 ;
    RECT -0.036 -0.028 0.036 0.028 ;
END V3_24x56_56V_56H

VIA V3_34x28_34V_28H
  LAYER m3 ;
    RECT -0.017 -0.038 0.017 0.038 ;
  LAYER v3 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER m4 ;
    RECT -0.041 -0.014 0.041 0.014 ;
END V3_34x28_34V_28H

VIA V3_34x28_44V_28H
  LAYER m3 ;
    RECT -0.022 -0.038 0.022 0.038 ;
  LAYER v3 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER m4 ;
    RECT -0.041 -0.014 0.041 0.014 ;
END V3_34x28_44V_28H

VIA V3_34x28_56H_28H
  LAYER m3 ;
    RECT -0.041 -0.028 0.041 0.028 ;
  LAYER v3 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER m4 ;
    RECT -0.041 -0.014 0.041 0.014 ;
END V3_34x28_56H_28H

VIA V3_34x28_56V_28H
  LAYER m3 ;
    RECT -0.028 -0.038 0.028 0.038 ;
  LAYER v3 ;
    RECT -0.017 -0.014 0.017 0.014 ;
  LAYER m4 ;
    RECT -0.041 -0.014 0.041 0.014 ;
END V3_34x28_56V_28H

VIA V3_35x35_44V_56H
  LAYER m3 ;
    RECT -0.022 -0.0415 0.022 0.0415 ;
  LAYER v3 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m4 ;
    RECT -0.0415 -0.028 0.0415 0.028 ;
END V3_35x35_44V_56H

VIA V3_35x35_44V_56V
  LAYER m3 ;
    RECT -0.022 -0.0415 0.022 0.0415 ;
  LAYER v3 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m4 ;
    RECT -0.028 -0.0415 0.028 0.0415 ;
END V3_35x35_44V_56V

VIA V3_35x35_56H_56H
  LAYER m3 ;
    RECT -0.0415 -0.028 0.0415 0.028 ;
  LAYER v3 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m4 ;
    RECT -0.0415 -0.028 0.0415 0.028 ;
END V3_35x35_56H_56H

VIA V3_35x35_56H_56V
  LAYER m3 ;
    RECT -0.0415 -0.028 0.0415 0.028 ;
  LAYER v3 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m4 ;
    RECT -0.028 -0.0415 0.028 0.0415 ;
END V3_35x35_56H_56V

VIA V3_35x35_56V_56H
  LAYER m3 ;
    RECT -0.028 -0.0415 0.028 0.0415 ;
  LAYER v3 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m4 ;
    RECT -0.0415 -0.028 0.0415 0.028 ;
END V3_35x35_56V_56H

VIA V3_35x35_56V_56V
  LAYER m3 ;
    RECT -0.028 -0.0415 0.028 0.0415 ;
  LAYER v3 ;
    RECT -0.0175 -0.0175 0.0175 0.0175 ;
  LAYER m4 ;
    RECT -0.028 -0.0415 0.028 0.0415 ;
END V3_35x35_56V_56V

VIA V4_120x24S_44H_120V
  LAYER m4 ;
    RECT -0.084 -0.022 0.084 0.022 ;
  LAYER v4 ;
    RECT -0.06 -0.012 0.06 0.012 ;
  LAYER m5 ;
    RECT -0.06 -0.05 0.06 0.05 ;
END V4_120x24S_44H_120V

VIA V4_120x24S_56H_120V
  LAYER m4 ;
    RECT -0.084 -0.028 0.084 0.028 ;
  LAYER v4 ;
    RECT -0.06 -0.012 0.06 0.012 ;
  LAYER m5 ;
    RECT -0.06 -0.05 0.06 0.05 ;
END V4_120x24S_56H_120V

VIA V4_120x24_44H_120H
  LAYER m4 ;
    RECT -0.084 -0.022 0.084 0.022 ;
  LAYER v4 ;
    RECT -0.06 -0.012 0.06 0.012 ;
  LAYER m5 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V4_120x24_44H_120H

VIA V4_120x24_44H_160H
  LAYER m4 ;
    RECT -0.084 -0.022 0.084 0.022 ;
  LAYER v4 ;
    RECT -0.06 -0.012 0.06 0.012 ;
  LAYER m5 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V4_120x24_44H_160H

VIA V4_120x24_44H_160V
  LAYER m4 ;
    RECT -0.084 -0.022 0.084 0.022 ;
  LAYER v4 ;
    RECT -0.06 -0.012 0.06 0.012 ;
  LAYER m5 ;
    RECT -0.08 -0.05 0.08 0.05 ;
END V4_120x24_44H_160V

VIA V4_120x24_44H_200H
  LAYER m4 ;
    RECT -0.084 -0.022 0.084 0.022 ;
  LAYER v4 ;
    RECT -0.06 -0.012 0.06 0.012 ;
  LAYER m5 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V4_120x24_44H_200H

VIA V4_120x24_44H_200V
  LAYER m4 ;
    RECT -0.084 -0.022 0.084 0.022 ;
  LAYER v4 ;
    RECT -0.06 -0.012 0.06 0.012 ;
  LAYER m5 ;
    RECT -0.1 -0.05 0.1 0.05 ;
END V4_120x24_44H_200V

VIA V4_120x24_44H_80H
  LAYER m4 ;
    RECT -0.084 -0.022 0.084 0.022 ;
  LAYER v4 ;
    RECT -0.06 -0.012 0.06 0.012 ;
  LAYER m5 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V4_120x24_44H_80H

VIA V4_120x24_56H_120H
  LAYER m4 ;
    RECT -0.084 -0.028 0.084 0.028 ;
  LAYER v4 ;
    RECT -0.06 -0.012 0.06 0.012 ;
  LAYER m5 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V4_120x24_56H_120H

VIA V4_120x24_56H_160H
  LAYER m4 ;
    RECT -0.084 -0.028 0.084 0.028 ;
  LAYER v4 ;
    RECT -0.06 -0.012 0.06 0.012 ;
  LAYER m5 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V4_120x24_56H_160H

VIA V4_120x24_56H_160V
  LAYER m4 ;
    RECT -0.084 -0.028 0.084 0.028 ;
  LAYER v4 ;
    RECT -0.06 -0.012 0.06 0.012 ;
  LAYER m5 ;
    RECT -0.08 -0.05 0.08 0.05 ;
END V4_120x24_56H_160V

VIA V4_120x24_56H_200H
  LAYER m4 ;
    RECT -0.084 -0.028 0.084 0.028 ;
  LAYER v4 ;
    RECT -0.06 -0.012 0.06 0.012 ;
  LAYER m5 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V4_120x24_56H_200H

VIA V4_120x24_56H_200V
  LAYER m4 ;
    RECT -0.084 -0.028 0.084 0.028 ;
  LAYER v4 ;
    RECT -0.06 -0.012 0.06 0.012 ;
  LAYER m5 ;
    RECT -0.1 -0.05 0.1 0.05 ;
END V4_120x24_56H_200V

VIA V4_120x24_56H_80H
  LAYER m4 ;
    RECT -0.084 -0.028 0.084 0.028 ;
  LAYER v4 ;
    RECT -0.06 -0.012 0.06 0.012 ;
  LAYER m5 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V4_120x24_56H_80H

VIA V4_40x24S_24H_40V
  LAYER m4 ;
    RECT -0.044 -0.012 0.044 0.012 ;
  LAYER v4 ;
    RECT -0.02 -0.012 0.02 0.012 ;
  LAYER m5 ;
    RECT -0.02 -0.05 0.02 0.05 ;
END V4_40x24S_24H_40V

VIA V4_40x24S_28H_40V
  LAYER m4 ;
    RECT -0.044 -0.014 0.044 0.014 ;
  LAYER v4 ;
    RECT -0.02 -0.012 0.02 0.012 ;
  LAYER m5 ;
    RECT -0.02 -0.05 0.02 0.05 ;
END V4_40x24S_28H_40V

VIA V4_40x24S_44H_40V
  LAYER m4 ;
    RECT -0.044 -0.022 0.044 0.022 ;
  LAYER v4 ;
    RECT -0.02 -0.012 0.02 0.012 ;
  LAYER m5 ;
    RECT -0.02 -0.05 0.02 0.05 ;
END V4_40x24S_44H_40V

VIA V4_40x24S_56H_40V
  LAYER m4 ;
    RECT -0.044 -0.028 0.044 0.028 ;
  LAYER v4 ;
    RECT -0.02 -0.012 0.02 0.012 ;
  LAYER m5 ;
    RECT -0.02 -0.05 0.02 0.05 ;
END V4_40x24S_56H_40V

VIA V4_40x24S_56V_40V
  LAYER m4 ;
    RECT -0.028 -0.036 0.028 0.036 ;
  LAYER v4 ;
    RECT -0.02 -0.012 0.02 0.012 ;
  LAYER m5 ;
    RECT -0.02 -0.05 0.02 0.05 ;
END V4_40x24S_56V_40V

VIA V4_40x28S_28H_40V
  LAYER m4 ;
    RECT -0.044 -0.014 0.044 0.014 ;
  LAYER v4 ;
    RECT -0.02 -0.014 0.02 0.014 ;
  LAYER m5 ;
    RECT -0.02 -0.052 0.02 0.052 ;
END V4_40x28S_28H_40V

VIA V4_40x28S_44H_40V
  LAYER m4 ;
    RECT -0.044 -0.022 0.044 0.022 ;
  LAYER v4 ;
    RECT -0.02 -0.014 0.02 0.014 ;
  LAYER m5 ;
    RECT -0.02 -0.052 0.02 0.052 ;
END V4_40x28S_44H_40V

VIA V4_40x28S_56H_40V
  LAYER m4 ;
    RECT -0.044 -0.028 0.044 0.028 ;
  LAYER v4 ;
    RECT -0.02 -0.014 0.02 0.014 ;
  LAYER m5 ;
    RECT -0.02 -0.052 0.02 0.052 ;
END V4_40x28S_56H_40V

VIA V4_40x28S_56V_40V
  LAYER m4 ;
    RECT -0.028 -0.038 0.028 0.038 ;
  LAYER v4 ;
    RECT -0.02 -0.014 0.02 0.014 ;
  LAYER m5 ;
    RECT -0.02 -0.052 0.02 0.052 ;
END V4_40x28S_56V_40V

VIA V4_60x24S_24H_60V
  LAYER m4 ;
    RECT -0.054 -0.012 0.054 0.012 ;
  LAYER v4 ;
    RECT -0.03 -0.012 0.03 0.012 ;
  LAYER m5 ;
    RECT -0.03 -0.05 0.03 0.05 ;
END V4_60x24S_24H_60V

VIA V4_60x24S_28H_60V
  LAYER m4 ;
    RECT -0.054 -0.014 0.054 0.014 ;
  LAYER v4 ;
    RECT -0.03 -0.012 0.03 0.012 ;
  LAYER m5 ;
    RECT -0.03 -0.05 0.03 0.05 ;
END V4_60x24S_28H_60V

VIA V4_60x24S_44H_60V
  LAYER m4 ;
    RECT -0.054 -0.022 0.054 0.022 ;
  LAYER v4 ;
    RECT -0.03 -0.012 0.03 0.012 ;
  LAYER m5 ;
    RECT -0.03 -0.05 0.03 0.05 ;
END V4_60x24S_44H_60V

VIA V4_60x24S_56H_60V
  LAYER m4 ;
    RECT -0.054 -0.028 0.054 0.028 ;
  LAYER v4 ;
    RECT -0.03 -0.012 0.03 0.012 ;
  LAYER m5 ;
    RECT -0.03 -0.05 0.03 0.05 ;
END V4_60x24S_56H_60V

VIA V4_80x24S_24H_80V
  LAYER m4 ;
    RECT -0.064 -0.012 0.064 0.012 ;
  LAYER v4 ;
    RECT -0.04 -0.012 0.04 0.012 ;
  LAYER m5 ;
    RECT -0.04 -0.05 0.04 0.05 ;
END V4_80x24S_24H_80V

VIA V4_80x24S_28H_80V
  LAYER m4 ;
    RECT -0.064 -0.014 0.064 0.014 ;
  LAYER v4 ;
    RECT -0.04 -0.012 0.04 0.012 ;
  LAYER m5 ;
    RECT -0.04 -0.05 0.04 0.05 ;
END V4_80x24S_28H_80V

VIA V4_80x24S_44H_80V
  LAYER m4 ;
    RECT -0.064 -0.022 0.064 0.022 ;
  LAYER v4 ;
    RECT -0.04 -0.012 0.04 0.012 ;
  LAYER m5 ;
    RECT -0.04 -0.05 0.04 0.05 ;
END V4_80x24S_44H_80V

VIA V4_80x24S_56H_80V
  LAYER m4 ;
    RECT -0.064 -0.028 0.064 0.028 ;
  LAYER v4 ;
    RECT -0.04 -0.012 0.04 0.012 ;
  LAYER m5 ;
    RECT -0.04 -0.05 0.04 0.05 ;
END V4_80x24S_56H_80V

VIA V5_120x40S_120H_120V
  LAYER m5 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V5_120x40S_120H_120V

VIA V5_120x40S_120V_120V
  LAYER m5 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V5_120x40S_120V_120V

VIA V5_120x40S_160H_120V
  LAYER m5 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V5_120x40S_160H_120V

VIA V5_120x40S_160V_120V
  LAYER m5 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V5_120x40S_160V_120V

VIA V5_120x40S_200H_120V
  LAYER m5 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V5_120x40S_200H_120V

VIA V5_120x40S_200V_120V
  LAYER m5 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V5_120x40S_200V_120V

VIA V5_120x40S_80H_120V
  LAYER m5 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V5_120x40S_80H_120V

VIA V5_120x40_120H_120H
  LAYER m5 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V5_120x40_120H_120H

VIA V5_120x40_120H_160H
  LAYER m5 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V5_120x40_120H_160H

VIA V5_120x40_120H_160V
  LAYER m5 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V5_120x40_120H_160V

VIA V5_120x40_120H_200H
  LAYER m5 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V5_120x40_120H_200H

VIA V5_120x40_120H_200V
  LAYER m5 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V5_120x40_120H_200V

VIA V5_120x40_120H_80H
  LAYER m5 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V5_120x40_120H_80H

VIA V5_120x40_160H_120H
  LAYER m5 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V5_120x40_160H_120H

VIA V5_120x40_160H_160H
  LAYER m5 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V5_120x40_160H_160H

VIA V5_120x40_160H_160V
  LAYER m5 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V5_120x40_160H_160V

VIA V5_120x40_160H_200H
  LAYER m5 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V5_120x40_160H_200H

VIA V5_120x40_160H_200V
  LAYER m5 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V5_120x40_160H_200V

VIA V5_120x40_160H_80H
  LAYER m5 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V5_120x40_160H_80H

VIA V5_120x40_160V_120H
  LAYER m5 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V5_120x40_160V_120H

VIA V5_120x40_160V_160H
  LAYER m5 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V5_120x40_160V_160H

VIA V5_120x40_160V_160V
  LAYER m5 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V5_120x40_160V_160V

VIA V5_120x40_160V_200H
  LAYER m5 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V5_120x40_160V_200H

VIA V5_120x40_160V_200V
  LAYER m5 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V5_120x40_160V_200V

VIA V5_120x40_160V_80H
  LAYER m5 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V5_120x40_160V_80H

VIA V5_120x40_200H_120H
  LAYER m5 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V5_120x40_200H_120H

VIA V5_120x40_200H_160H
  LAYER m5 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V5_120x40_200H_160H

VIA V5_120x40_200H_160V
  LAYER m5 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V5_120x40_200H_160V

VIA V5_120x40_200H_200H
  LAYER m5 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V5_120x40_200H_200H

VIA V5_120x40_200H_200V
  LAYER m5 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V5_120x40_200H_200V

VIA V5_120x40_200H_80H
  LAYER m5 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V5_120x40_200H_80H

VIA V5_120x40_200V_120H
  LAYER m5 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V5_120x40_200V_120H

VIA V5_120x40_200V_160H
  LAYER m5 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V5_120x40_200V_160H

VIA V5_120x40_200V_160V
  LAYER m5 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V5_120x40_200V_160V

VIA V5_120x40_200V_200H
  LAYER m5 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V5_120x40_200V_200H

VIA V5_120x40_200V_200V
  LAYER m5 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V5_120x40_200V_200V

VIA V5_120x40_200V_80H
  LAYER m5 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V5_120x40_200V_80H

VIA V5_120x40_80H_120H
  LAYER m5 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V5_120x40_80H_120H

VIA V5_120x40_80H_160H
  LAYER m5 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V5_120x40_80H_160H

VIA V5_120x40_80H_160V
  LAYER m5 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V5_120x40_80H_160V

VIA V5_120x40_80H_200H
  LAYER m5 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V5_120x40_80H_200H

VIA V5_120x40_80H_200V
  LAYER m5 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V5_120x40_80H_200V

VIA V5_120x40_80H_80H
  LAYER m5 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v5 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m6 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V5_120x40_80H_80H

VIA V5_40Sx120_120H_120H
  LAYER m5 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V5_40Sx120_120H_120H

VIA V5_40Sx120_120V_120H
  LAYER m5 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V5_40Sx120_120V_120H

VIA V5_40Sx120_160H_120H
  LAYER m5 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V5_40Sx120_160H_120H

VIA V5_40Sx120_160V_120H
  LAYER m5 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V5_40Sx120_160V_120H

VIA V5_40Sx120_200H_120H
  LAYER m5 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V5_40Sx120_200H_120H

VIA V5_40Sx120_200V_120H
  LAYER m5 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V5_40Sx120_200V_120H

VIA V5_40Sx120_40V_120H
  LAYER m5 ;
    RECT -0.02 -0.084 0.02 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V5_40Sx120_40V_120H

VIA V5_40Sx120_60V_120H
  LAYER m5 ;
    RECT -0.03 -0.084 0.03 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V5_40Sx120_60V_120H

VIA V5_40Sx120_80V_120H
  LAYER m5 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V5_40Sx120_80V_120H

VIA V5_40Sx40_120H_40H
  LAYER m5 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v5 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m6 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V5_40Sx40_120H_40H

VIA V5_40Sx40_120V_40H
  LAYER m5 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v5 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m6 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V5_40Sx40_120V_40H

VIA V5_40Sx40_160H_40H
  LAYER m5 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v5 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m6 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V5_40Sx40_160H_40H

VIA V5_40Sx40_160V_40H
  LAYER m5 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v5 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m6 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V5_40Sx40_160V_40H

VIA V5_40Sx40_200H_40H
  LAYER m5 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v5 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m6 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V5_40Sx40_200H_40H

VIA V5_40Sx40_200V_40H
  LAYER m5 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v5 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m6 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V5_40Sx40_200V_40H

VIA V5_40Sx40_40V_40H
  LAYER m5 ;
    RECT -0.02 -0.044 0.02 0.044 ;
  LAYER v5 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m6 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V5_40Sx40_40V_40H

VIA V5_40Sx40_60V_40H
  LAYER m5 ;
    RECT -0.03 -0.044 0.03 0.044 ;
  LAYER v5 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m6 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V5_40Sx40_60V_40H

VIA V5_40Sx40_80H_40H
  LAYER m5 ;
    RECT -0.044 -0.04 0.044 0.04 ;
  LAYER v5 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m6 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V5_40Sx40_80H_40H

VIA V5_40Sx40_80V_40H
  LAYER m5 ;
    RECT -0.04 -0.044 0.04 0.044 ;
  LAYER v5 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m6 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V5_40Sx40_80V_40H

VIA V5_40Sx60_120H_60H
  LAYER m5 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v5 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m6 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V5_40Sx60_120H_60H

VIA V5_40Sx60_120V_60H
  LAYER m5 ;
    RECT -0.06 -0.054 0.06 0.054 ;
  LAYER v5 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m6 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V5_40Sx60_120V_60H

VIA V5_40Sx60_160H_60H
  LAYER m5 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v5 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m6 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V5_40Sx60_160H_60H

VIA V5_40Sx60_160V_60H
  LAYER m5 ;
    RECT -0.08 -0.054 0.08 0.054 ;
  LAYER v5 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m6 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V5_40Sx60_160V_60H

VIA V5_40Sx60_200H_60H
  LAYER m5 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v5 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m6 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V5_40Sx60_200H_60H

VIA V5_40Sx60_200V_60H
  LAYER m5 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v5 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m6 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V5_40Sx60_200V_60H

VIA V5_40Sx60_40V_60H
  LAYER m5 ;
    RECT -0.02 -0.054 0.02 0.054 ;
  LAYER v5 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m6 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V5_40Sx60_40V_60H

VIA V5_40Sx60_60V_60H
  LAYER m5 ;
    RECT -0.03 -0.054 0.03 0.054 ;
  LAYER v5 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m6 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V5_40Sx60_60V_60H

VIA V5_40Sx60_80H_60H
  LAYER m5 ;
    RECT -0.044 -0.04 0.044 0.04 ;
  LAYER v5 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m6 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V5_40Sx60_80H_60H

VIA V5_40Sx60_80V_60H
  LAYER m5 ;
    RECT -0.04 -0.054 0.04 0.054 ;
  LAYER v5 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m6 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V5_40Sx60_80V_60H

VIA V5_40Sx80_120H_80H
  LAYER m5 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v5 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m6 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V5_40Sx80_120H_80H

VIA V5_40Sx80_120V_80H
  LAYER m5 ;
    RECT -0.06 -0.064 0.06 0.064 ;
  LAYER v5 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m6 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V5_40Sx80_120V_80H

VIA V5_40Sx80_160H_80H
  LAYER m5 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v5 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m6 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V5_40Sx80_160H_80H

VIA V5_40Sx80_160V_80H
  LAYER m5 ;
    RECT -0.08 -0.064 0.08 0.064 ;
  LAYER v5 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m6 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V5_40Sx80_160V_80H

VIA V5_40Sx80_200H_80H
  LAYER m5 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v5 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m6 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V5_40Sx80_200H_80H

VIA V5_40Sx80_200V_80H
  LAYER m5 ;
    RECT -0.1 -0.064 0.1 0.064 ;
  LAYER v5 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m6 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V5_40Sx80_200V_80H

VIA V5_40Sx80_40V_80H
  LAYER m5 ;
    RECT -0.02 -0.064 0.02 0.064 ;
  LAYER v5 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m6 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V5_40Sx80_40V_80H

VIA V5_40Sx80_60V_80H
  LAYER m5 ;
    RECT -0.03 -0.064 0.03 0.064 ;
  LAYER v5 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m6 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V5_40Sx80_60V_80H

VIA V5_40Sx80_80H_80H
  LAYER m5 ;
    RECT -0.044 -0.04 0.044 0.04 ;
  LAYER v5 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m6 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V5_40Sx80_80H_80H

VIA V5_40Sx80_80V_80H
  LAYER m5 ;
    RECT -0.04 -0.064 0.04 0.064 ;
  LAYER v5 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m6 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V5_40Sx80_80V_80H

VIA V5_40x120_120V_120V
  LAYER m5 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V5_40x120_120V_120V

VIA V5_40x120_120V_160H
  LAYER m5 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V5_40x120_120V_160H

VIA V5_40x120_120V_160V
  LAYER m5 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V5_40x120_120V_160V

VIA V5_40x120_120V_200H
  LAYER m5 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V5_40x120_120V_200H

VIA V5_40x120_120V_200V
  LAYER m5 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V5_40x120_120V_200V

VIA V5_40x120_120V_80V
  LAYER m5 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V5_40x120_120V_80V

VIA V5_40x120_160H_120V
  LAYER m5 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V5_40x120_160H_120V

VIA V5_40x120_160H_160H
  LAYER m5 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V5_40x120_160H_160H

VIA V5_40x120_160H_160V
  LAYER m5 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V5_40x120_160H_160V

VIA V5_40x120_160H_200H
  LAYER m5 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V5_40x120_160H_200H

VIA V5_40x120_160H_200V
  LAYER m5 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V5_40x120_160H_200V

VIA V5_40x120_160H_80V
  LAYER m5 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V5_40x120_160H_80V

VIA V5_40x120_160V_120V
  LAYER m5 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V5_40x120_160V_120V

VIA V5_40x120_160V_160H
  LAYER m5 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V5_40x120_160V_160H

VIA V5_40x120_160V_160V
  LAYER m5 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V5_40x120_160V_160V

VIA V5_40x120_160V_200H
  LAYER m5 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V5_40x120_160V_200H

VIA V5_40x120_160V_200V
  LAYER m5 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V5_40x120_160V_200V

VIA V5_40x120_160V_80V
  LAYER m5 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V5_40x120_160V_80V

VIA V5_40x120_200H_120V
  LAYER m5 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V5_40x120_200H_120V

VIA V5_40x120_200H_160H
  LAYER m5 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V5_40x120_200H_160H

VIA V5_40x120_200H_160V
  LAYER m5 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V5_40x120_200H_160V

VIA V5_40x120_200H_200H
  LAYER m5 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V5_40x120_200H_200H

VIA V5_40x120_200H_200V
  LAYER m5 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V5_40x120_200H_200V

VIA V5_40x120_200H_80V
  LAYER m5 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V5_40x120_200H_80V

VIA V5_40x120_200V_120V
  LAYER m5 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V5_40x120_200V_120V

VIA V5_40x120_200V_160H
  LAYER m5 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V5_40x120_200V_160H

VIA V5_40x120_200V_160V
  LAYER m5 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V5_40x120_200V_160V

VIA V5_40x120_200V_200H
  LAYER m5 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V5_40x120_200V_200H

VIA V5_40x120_200V_200V
  LAYER m5 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V5_40x120_200V_200V

VIA V5_40x120_200V_80V
  LAYER m5 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V5_40x120_200V_80V

VIA V5_40x120_80V_120V
  LAYER m5 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V5_40x120_80V_120V

VIA V5_40x120_80V_160H
  LAYER m5 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V5_40x120_80V_160H

VIA V5_40x120_80V_160V
  LAYER m5 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V5_40x120_80V_160V

VIA V5_40x120_80V_200H
  LAYER m5 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V5_40x120_80V_200H

VIA V5_40x120_80V_200V
  LAYER m5 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V5_40x120_80V_200V

VIA V5_40x120_80V_80V
  LAYER m5 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v5 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m6 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V5_40x120_80V_80V

VIA V5_60Sx40_120H_40H
  LAYER m5 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v5 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m6 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V5_60Sx40_120H_40H

VIA V5_60Sx40_120V_40H
  LAYER m5 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v5 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m6 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V5_60Sx40_120V_40H

VIA V5_60Sx40_160H_40H
  LAYER m5 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v5 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m6 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V5_60Sx40_160H_40H

VIA V5_60Sx40_160V_40H
  LAYER m5 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v5 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m6 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V5_60Sx40_160V_40H

VIA V5_60Sx40_200H_40H
  LAYER m5 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v5 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m6 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V5_60Sx40_200H_40H

VIA V5_60Sx40_200V_40H
  LAYER m5 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v5 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m6 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V5_60Sx40_200V_40H

VIA V5_60Sx40_60V_40H
  LAYER m5 ;
    RECT -0.03 -0.044 0.03 0.044 ;
  LAYER v5 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m6 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V5_60Sx40_60V_40H

VIA V5_60Sx40_80H_40H
  LAYER m5 ;
    RECT -0.054 -0.04 0.054 0.04 ;
  LAYER v5 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m6 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V5_60Sx40_80H_40H

VIA V5_60Sx40_80V_40H
  LAYER m5 ;
    RECT -0.04 -0.044 0.04 0.044 ;
  LAYER v5 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m6 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V5_60Sx40_80V_40H

VIA V5_60Sx60_120H_60H
  LAYER m5 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v5 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m6 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V5_60Sx60_120H_60H

VIA V5_60Sx60_120V_60H
  LAYER m5 ;
    RECT -0.06 -0.054 0.06 0.054 ;
  LAYER v5 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m6 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V5_60Sx60_120V_60H

VIA V5_60Sx60_160H_60H
  LAYER m5 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v5 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m6 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V5_60Sx60_160H_60H

VIA V5_60Sx60_160V_60H
  LAYER m5 ;
    RECT -0.08 -0.054 0.08 0.054 ;
  LAYER v5 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m6 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V5_60Sx60_160V_60H

VIA V5_60Sx60_200H_60H
  LAYER m5 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v5 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m6 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V5_60Sx60_200H_60H

VIA V5_60Sx60_200V_60H
  LAYER m5 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v5 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m6 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V5_60Sx60_200V_60H

VIA V5_60Sx60_60V_60H
  LAYER m5 ;
    RECT -0.03 -0.054 0.03 0.054 ;
  LAYER v5 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m6 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V5_60Sx60_60V_60H

VIA V5_60Sx60_80H_60H
  LAYER m5 ;
    RECT -0.054 -0.04 0.054 0.04 ;
  LAYER v5 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m6 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V5_60Sx60_80H_60H

VIA V5_60Sx60_80V_60H
  LAYER m5 ;
    RECT -0.04 -0.054 0.04 0.054 ;
  LAYER v5 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m6 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V5_60Sx60_80V_60H

VIA V5_60Sx80_120H_80H
  LAYER m5 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v5 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m6 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V5_60Sx80_120H_80H

VIA V5_60Sx80_120V_80H
  LAYER m5 ;
    RECT -0.06 -0.064 0.06 0.064 ;
  LAYER v5 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m6 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V5_60Sx80_120V_80H

VIA V5_60Sx80_160H_80H
  LAYER m5 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v5 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m6 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V5_60Sx80_160H_80H

VIA V5_60Sx80_160V_80H
  LAYER m5 ;
    RECT -0.08 -0.064 0.08 0.064 ;
  LAYER v5 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m6 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V5_60Sx80_160V_80H

VIA V5_60Sx80_200H_80H
  LAYER m5 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v5 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m6 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V5_60Sx80_200H_80H

VIA V5_60Sx80_200V_80H
  LAYER m5 ;
    RECT -0.1 -0.064 0.1 0.064 ;
  LAYER v5 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m6 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V5_60Sx80_200V_80H

VIA V5_60Sx80_60V_80H
  LAYER m5 ;
    RECT -0.03 -0.064 0.03 0.064 ;
  LAYER v5 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m6 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V5_60Sx80_60V_80H

VIA V5_60Sx80_80H_80H
  LAYER m5 ;
    RECT -0.054 -0.04 0.054 0.04 ;
  LAYER v5 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m6 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V5_60Sx80_80H_80H

VIA V5_60Sx80_80V_80H
  LAYER m5 ;
    RECT -0.04 -0.064 0.04 0.064 ;
  LAYER v5 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m6 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V5_60Sx80_80V_80H

VIA V5_80x40S_120H_80V
  LAYER m5 ;
    RECT -0.064 -0.06 0.064 0.06 ;
  LAYER v5 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m6 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V5_80x40S_120H_80V

VIA V5_80x40S_120V_80V
  LAYER m5 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v5 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m6 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V5_80x40S_120V_80V

VIA V5_80x40S_160H_80V
  LAYER m5 ;
    RECT -0.064 -0.08 0.064 0.08 ;
  LAYER v5 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m6 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V5_80x40S_160H_80V

VIA V5_80x40S_160V_80V
  LAYER m5 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v5 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m6 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V5_80x40S_160V_80V

VIA V5_80x40S_200H_80V
  LAYER m5 ;
    RECT -0.064 -0.1 0.064 0.1 ;
  LAYER v5 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m6 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V5_80x40S_200H_80V

VIA V5_80x40S_200V_80V
  LAYER m5 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v5 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m6 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V5_80x40S_200V_80V

VIA V5_80x40S_80H_80V
  LAYER m5 ;
    RECT -0.064 -0.04 0.064 0.04 ;
  LAYER v5 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m6 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V5_80x40S_80H_80V

VIA V5_80x40S_80V_80V
  LAYER m5 ;
    RECT -0.04 -0.044 0.04 0.044 ;
  LAYER v5 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m6 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V5_80x40S_80V_80V

VIA V6_120x40S_120H_120V
  LAYER m6 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V6_120x40S_120H_120V

VIA V6_120x40S_120V_120V
  LAYER m6 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V6_120x40S_120V_120V

VIA V6_120x40S_160H_120V
  LAYER m6 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V6_120x40S_160H_120V

VIA V6_120x40S_160V_120V
  LAYER m6 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V6_120x40S_160V_120V

VIA V6_120x40S_200H_120V
  LAYER m6 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V6_120x40S_200H_120V

VIA V6_120x40S_200V_120V
  LAYER m6 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V6_120x40S_200V_120V

VIA V6_120x40S_40H_120V
  LAYER m6 ;
    RECT -0.084 -0.02 0.084 0.02 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V6_120x40S_40H_120V

VIA V6_120x40S_60H_120V
  LAYER m6 ;
    RECT -0.084 -0.03 0.084 0.03 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V6_120x40S_60H_120V

VIA V6_120x40S_80H_120V
  LAYER m6 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V6_120x40S_80H_120V

VIA V6_120x40_120H_120H
  LAYER m6 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V6_120x40_120H_120H

VIA V6_120x40_120H_160H
  LAYER m6 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V6_120x40_120H_160H

VIA V6_120x40_120H_160V
  LAYER m6 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V6_120x40_120H_160V

VIA V6_120x40_120H_200H
  LAYER m6 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V6_120x40_120H_200H

VIA V6_120x40_120H_200V
  LAYER m6 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V6_120x40_120H_200V

VIA V6_120x40_120H_80H
  LAYER m6 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V6_120x40_120H_80H

VIA V6_120x40_160H_120H
  LAYER m6 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V6_120x40_160H_120H

VIA V6_120x40_160H_160H
  LAYER m6 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V6_120x40_160H_160H

VIA V6_120x40_160H_160V
  LAYER m6 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V6_120x40_160H_160V

VIA V6_120x40_160H_200H
  LAYER m6 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V6_120x40_160H_200H

VIA V6_120x40_160H_200V
  LAYER m6 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V6_120x40_160H_200V

VIA V6_120x40_160H_80H
  LAYER m6 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V6_120x40_160H_80H

VIA V6_120x40_160V_120H
  LAYER m6 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V6_120x40_160V_120H

VIA V6_120x40_160V_160H
  LAYER m6 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V6_120x40_160V_160H

VIA V6_120x40_160V_160V
  LAYER m6 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V6_120x40_160V_160V

VIA V6_120x40_160V_200H
  LAYER m6 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V6_120x40_160V_200H

VIA V6_120x40_160V_200V
  LAYER m6 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V6_120x40_160V_200V

VIA V6_120x40_160V_80H
  LAYER m6 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V6_120x40_160V_80H

VIA V6_120x40_200H_120H
  LAYER m6 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V6_120x40_200H_120H

VIA V6_120x40_200H_160H
  LAYER m6 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V6_120x40_200H_160H

VIA V6_120x40_200H_160V
  LAYER m6 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V6_120x40_200H_160V

VIA V6_120x40_200H_200H
  LAYER m6 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V6_120x40_200H_200H

VIA V6_120x40_200H_200V
  LAYER m6 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V6_120x40_200H_200V

VIA V6_120x40_200H_80H
  LAYER m6 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V6_120x40_200H_80H

VIA V6_120x40_200V_120H
  LAYER m6 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V6_120x40_200V_120H

VIA V6_120x40_200V_160H
  LAYER m6 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V6_120x40_200V_160H

VIA V6_120x40_200V_160V
  LAYER m6 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V6_120x40_200V_160V

VIA V6_120x40_200V_200H
  LAYER m6 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V6_120x40_200V_200H

VIA V6_120x40_200V_200V
  LAYER m6 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V6_120x40_200V_200V

VIA V6_120x40_200V_80H
  LAYER m6 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V6_120x40_200V_80H

VIA V6_120x40_80H_120H
  LAYER m6 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V6_120x40_80H_120H

VIA V6_120x40_80H_160H
  LAYER m6 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V6_120x40_80H_160H

VIA V6_120x40_80H_160V
  LAYER m6 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V6_120x40_80H_160V

VIA V6_120x40_80H_200H
  LAYER m6 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V6_120x40_80H_200H

VIA V6_120x40_80H_200V
  LAYER m6 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V6_120x40_80H_200V

VIA V6_120x40_80H_80H
  LAYER m6 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v6 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m7 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V6_120x40_80H_80H

VIA V6_40Sx120_120H_120H
  LAYER m6 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V6_40Sx120_120H_120H

VIA V6_40Sx120_120V_120H
  LAYER m6 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V6_40Sx120_120V_120H

VIA V6_40Sx120_160H_120H
  LAYER m6 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V6_40Sx120_160H_120H

VIA V6_40Sx120_160V_120H
  LAYER m6 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V6_40Sx120_160V_120H

VIA V6_40Sx120_200H_120H
  LAYER m6 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V6_40Sx120_200H_120H

VIA V6_40Sx120_200V_120H
  LAYER m6 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V6_40Sx120_200V_120H

VIA V6_40Sx120_80V_120H
  LAYER m6 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V6_40Sx120_80V_120H

VIA V6_40Sx80_120H_80H
  LAYER m6 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v6 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m7 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V6_40Sx80_120H_80H

VIA V6_40Sx80_120V_80H
  LAYER m6 ;
    RECT -0.06 -0.064 0.06 0.064 ;
  LAYER v6 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m7 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V6_40Sx80_120V_80H

VIA V6_40Sx80_160H_80H
  LAYER m6 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v6 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m7 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V6_40Sx80_160H_80H

VIA V6_40Sx80_160V_80H
  LAYER m6 ;
    RECT -0.08 -0.064 0.08 0.064 ;
  LAYER v6 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m7 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V6_40Sx80_160V_80H

VIA V6_40Sx80_200H_80H
  LAYER m6 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v6 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m7 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V6_40Sx80_200H_80H

VIA V6_40Sx80_200V_80H
  LAYER m6 ;
    RECT -0.1 -0.064 0.1 0.064 ;
  LAYER v6 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m7 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V6_40Sx80_200V_80H

VIA V6_40Sx80_80H_80H
  LAYER m6 ;
    RECT -0.044 -0.04 0.044 0.04 ;
  LAYER v6 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m7 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V6_40Sx80_80H_80H

VIA V6_40Sx80_80V_80H
  LAYER m6 ;
    RECT -0.04 -0.064 0.04 0.064 ;
  LAYER v6 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m7 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V6_40Sx80_80V_80H

VIA V6_40x120_120V_120V
  LAYER m6 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V6_40x120_120V_120V

VIA V6_40x120_120V_160H
  LAYER m6 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V6_40x120_120V_160H

VIA V6_40x120_120V_160V
  LAYER m6 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V6_40x120_120V_160V

VIA V6_40x120_120V_200H
  LAYER m6 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V6_40x120_120V_200H

VIA V6_40x120_120V_200V
  LAYER m6 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V6_40x120_120V_200V

VIA V6_40x120_120V_80V
  LAYER m6 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V6_40x120_120V_80V

VIA V6_40x120_160H_120V
  LAYER m6 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V6_40x120_160H_120V

VIA V6_40x120_160H_160H
  LAYER m6 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V6_40x120_160H_160H

VIA V6_40x120_160H_160V
  LAYER m6 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V6_40x120_160H_160V

VIA V6_40x120_160H_200H
  LAYER m6 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V6_40x120_160H_200H

VIA V6_40x120_160H_200V
  LAYER m6 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V6_40x120_160H_200V

VIA V6_40x120_160H_80V
  LAYER m6 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V6_40x120_160H_80V

VIA V6_40x120_160V_120V
  LAYER m6 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V6_40x120_160V_120V

VIA V6_40x120_160V_160H
  LAYER m6 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V6_40x120_160V_160H

VIA V6_40x120_160V_160V
  LAYER m6 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V6_40x120_160V_160V

VIA V6_40x120_160V_200H
  LAYER m6 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V6_40x120_160V_200H

VIA V6_40x120_160V_200V
  LAYER m6 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V6_40x120_160V_200V

VIA V6_40x120_160V_80V
  LAYER m6 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V6_40x120_160V_80V

VIA V6_40x120_200H_120V
  LAYER m6 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V6_40x120_200H_120V

VIA V6_40x120_200H_160H
  LAYER m6 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V6_40x120_200H_160H

VIA V6_40x120_200H_160V
  LAYER m6 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V6_40x120_200H_160V

VIA V6_40x120_200H_200H
  LAYER m6 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V6_40x120_200H_200H

VIA V6_40x120_200H_200V
  LAYER m6 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V6_40x120_200H_200V

VIA V6_40x120_200H_80V
  LAYER m6 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V6_40x120_200H_80V

VIA V6_40x120_200V_120V
  LAYER m6 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V6_40x120_200V_120V

VIA V6_40x120_200V_160H
  LAYER m6 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V6_40x120_200V_160H

VIA V6_40x120_200V_160V
  LAYER m6 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V6_40x120_200V_160V

VIA V6_40x120_200V_200H
  LAYER m6 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V6_40x120_200V_200H

VIA V6_40x120_200V_200V
  LAYER m6 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V6_40x120_200V_200V

VIA V6_40x120_200V_80V
  LAYER m6 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V6_40x120_200V_80V

VIA V6_40x120_80V_120V
  LAYER m6 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V6_40x120_80V_120V

VIA V6_40x120_80V_160H
  LAYER m6 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V6_40x120_80V_160H

VIA V6_40x120_80V_160V
  LAYER m6 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V6_40x120_80V_160V

VIA V6_40x120_80V_200H
  LAYER m6 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V6_40x120_80V_200H

VIA V6_40x120_80V_200V
  LAYER m6 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V6_40x120_80V_200V

VIA V6_40x120_80V_80V
  LAYER m6 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v6 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m7 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V6_40x120_80V_80V

VIA V6_40x40S_120H_40V
  LAYER m6 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v6 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m7 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V6_40x40S_120H_40V

VIA V6_40x40S_120V_40V
  LAYER m6 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v6 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m7 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V6_40x40S_120V_40V

VIA V6_40x40S_160H_40V
  LAYER m6 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v6 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m7 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V6_40x40S_160H_40V

VIA V6_40x40S_160V_40V
  LAYER m6 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v6 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m7 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V6_40x40S_160V_40V

VIA V6_40x40S_200H_40V
  LAYER m6 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v6 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m7 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V6_40x40S_200H_40V

VIA V6_40x40S_200V_40V
  LAYER m6 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v6 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m7 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V6_40x40S_200V_40V

VIA V6_40x40S_40H_40V
  LAYER m6 ;
    RECT -0.044 -0.02 0.044 0.02 ;
  LAYER v6 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m7 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V6_40x40S_40H_40V

VIA V6_40x40S_60H_40V
  LAYER m6 ;
    RECT -0.044 -0.03 0.044 0.03 ;
  LAYER v6 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m7 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V6_40x40S_60H_40V

VIA V6_40x40S_80H_40V
  LAYER m6 ;
    RECT -0.044 -0.04 0.044 0.04 ;
  LAYER v6 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m7 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V6_40x40S_80H_40V

VIA V6_40x40S_80V_40V
  LAYER m6 ;
    RECT -0.04 -0.044 0.04 0.044 ;
  LAYER v6 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m7 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V6_40x40S_80V_40V

VIA V6_40x60S_120H_40V
  LAYER m6 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v6 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m7 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V6_40x60S_120H_40V

VIA V6_40x60S_120V_40V
  LAYER m6 ;
    RECT -0.06 -0.054 0.06 0.054 ;
  LAYER v6 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m7 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V6_40x60S_120V_40V

VIA V6_40x60S_160H_40V
  LAYER m6 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v6 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m7 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V6_40x60S_160H_40V

VIA V6_40x60S_160V_40V
  LAYER m6 ;
    RECT -0.08 -0.054 0.08 0.054 ;
  LAYER v6 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m7 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V6_40x60S_160V_40V

VIA V6_40x60S_200H_40V
  LAYER m6 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v6 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m7 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V6_40x60S_200H_40V

VIA V6_40x60S_200V_40V
  LAYER m6 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v6 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m7 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V6_40x60S_200V_40V

VIA V6_40x60S_60H_40V
  LAYER m6 ;
    RECT -0.044 -0.03 0.044 0.03 ;
  LAYER v6 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m7 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V6_40x60S_60H_40V

VIA V6_40x60S_80H_40V
  LAYER m6 ;
    RECT -0.044 -0.04 0.044 0.04 ;
  LAYER v6 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m7 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V6_40x60S_80H_40V

VIA V6_40x60S_80V_40V
  LAYER m6 ;
    RECT -0.04 -0.054 0.04 0.054 ;
  LAYER v6 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m7 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V6_40x60S_80V_40V

VIA V6_60x40S_120H_60V
  LAYER m6 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v6 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m7 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V6_60x40S_120H_60V

VIA V6_60x40S_120V_60V
  LAYER m6 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v6 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m7 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V6_60x40S_120V_60V

VIA V6_60x40S_160H_60V
  LAYER m6 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v6 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m7 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V6_60x40S_160H_60V

VIA V6_60x40S_160V_60V
  LAYER m6 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v6 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m7 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V6_60x40S_160V_60V

VIA V6_60x40S_200H_60V
  LAYER m6 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v6 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m7 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V6_60x40S_200H_60V

VIA V6_60x40S_200V_60V
  LAYER m6 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v6 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m7 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V6_60x40S_200V_60V

VIA V6_60x40S_40H_60V
  LAYER m6 ;
    RECT -0.054 -0.02 0.054 0.02 ;
  LAYER v6 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m7 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V6_60x40S_40H_60V

VIA V6_60x40S_60H_60V
  LAYER m6 ;
    RECT -0.054 -0.03 0.054 0.03 ;
  LAYER v6 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m7 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V6_60x40S_60H_60V

VIA V6_60x40S_80H_60V
  LAYER m6 ;
    RECT -0.054 -0.04 0.054 0.04 ;
  LAYER v6 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m7 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V6_60x40S_80H_60V

VIA V6_60x40S_80V_60V
  LAYER m6 ;
    RECT -0.04 -0.044 0.04 0.044 ;
  LAYER v6 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m7 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V6_60x40S_80V_60V

VIA V6_60x60S_120H_60V
  LAYER m6 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v6 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m7 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V6_60x60S_120H_60V

VIA V6_60x60S_120V_60V
  LAYER m6 ;
    RECT -0.06 -0.054 0.06 0.054 ;
  LAYER v6 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m7 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V6_60x60S_120V_60V

VIA V6_60x60S_160H_60V
  LAYER m6 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v6 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m7 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V6_60x60S_160H_60V

VIA V6_60x60S_160V_60V
  LAYER m6 ;
    RECT -0.08 -0.054 0.08 0.054 ;
  LAYER v6 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m7 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V6_60x60S_160V_60V

VIA V6_60x60S_200H_60V
  LAYER m6 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v6 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m7 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V6_60x60S_200H_60V

VIA V6_60x60S_200V_60V
  LAYER m6 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v6 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m7 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V6_60x60S_200V_60V

VIA V6_60x60S_60H_60V
  LAYER m6 ;
    RECT -0.054 -0.03 0.054 0.03 ;
  LAYER v6 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m7 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V6_60x60S_60H_60V

VIA V6_60x60S_80H_60V
  LAYER m6 ;
    RECT -0.054 -0.04 0.054 0.04 ;
  LAYER v6 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m7 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V6_60x60S_80H_60V

VIA V6_60x60S_80V_60V
  LAYER m6 ;
    RECT -0.04 -0.054 0.04 0.054 ;
  LAYER v6 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m7 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V6_60x60S_80V_60V

VIA V6_80x40S_120H_80V
  LAYER m6 ;
    RECT -0.064 -0.06 0.064 0.06 ;
  LAYER v6 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m7 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V6_80x40S_120H_80V

VIA V6_80x40S_120V_80V
  LAYER m6 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v6 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m7 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V6_80x40S_120V_80V

VIA V6_80x40S_160H_80V
  LAYER m6 ;
    RECT -0.064 -0.08 0.064 0.08 ;
  LAYER v6 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m7 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V6_80x40S_160H_80V

VIA V6_80x40S_160V_80V
  LAYER m6 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v6 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m7 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V6_80x40S_160V_80V

VIA V6_80x40S_200H_80V
  LAYER m6 ;
    RECT -0.064 -0.1 0.064 0.1 ;
  LAYER v6 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m7 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V6_80x40S_200H_80V

VIA V6_80x40S_200V_80V
  LAYER m6 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v6 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m7 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V6_80x40S_200V_80V

VIA V6_80x40S_40H_80V
  LAYER m6 ;
    RECT -0.064 -0.02 0.064 0.02 ;
  LAYER v6 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m7 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V6_80x40S_40H_80V

VIA V6_80x40S_60H_80V
  LAYER m6 ;
    RECT -0.064 -0.03 0.064 0.03 ;
  LAYER v6 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m7 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V6_80x40S_60H_80V

VIA V6_80x40S_80H_80V
  LAYER m6 ;
    RECT -0.064 -0.04 0.064 0.04 ;
  LAYER v6 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m7 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V6_80x40S_80H_80V

VIA V6_80x40S_80V_80V
  LAYER m6 ;
    RECT -0.04 -0.044 0.04 0.044 ;
  LAYER v6 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m7 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V6_80x40S_80V_80V

VIA V6_80x60S_120H_80V
  LAYER m6 ;
    RECT -0.064 -0.06 0.064 0.06 ;
  LAYER v6 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m7 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V6_80x60S_120H_80V

VIA V6_80x60S_120V_80V
  LAYER m6 ;
    RECT -0.06 -0.054 0.06 0.054 ;
  LAYER v6 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m7 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V6_80x60S_120V_80V

VIA V6_80x60S_160H_80V
  LAYER m6 ;
    RECT -0.064 -0.08 0.064 0.08 ;
  LAYER v6 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m7 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V6_80x60S_160H_80V

VIA V6_80x60S_160V_80V
  LAYER m6 ;
    RECT -0.08 -0.054 0.08 0.054 ;
  LAYER v6 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m7 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V6_80x60S_160V_80V

VIA V6_80x60S_200H_80V
  LAYER m6 ;
    RECT -0.064 -0.1 0.064 0.1 ;
  LAYER v6 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m7 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V6_80x60S_200H_80V

VIA V6_80x60S_200V_80V
  LAYER m6 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v6 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m7 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V6_80x60S_200V_80V

VIA V6_80x60S_60H_80V
  LAYER m6 ;
    RECT -0.064 -0.03 0.064 0.03 ;
  LAYER v6 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m7 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V6_80x60S_60H_80V

VIA V6_80x60S_80H_80V
  LAYER m6 ;
    RECT -0.064 -0.04 0.064 0.04 ;
  LAYER v6 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m7 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V6_80x60S_80H_80V

VIA V6_80x60S_80V_80V
  LAYER m6 ;
    RECT -0.04 -0.054 0.04 0.054 ;
  LAYER v6 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m7 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V6_80x60S_80V_80V

VIA V7_120x40S_120H_120V
  LAYER m7 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V7_120x40S_120H_120V

VIA V7_120x40S_120V_120V
  LAYER m7 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V7_120x40S_120V_120V

VIA V7_120x40S_160H_120V
  LAYER m7 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V7_120x40S_160H_120V

VIA V7_120x40S_160V_120V
  LAYER m7 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V7_120x40S_160V_120V

VIA V7_120x40S_200H_120V
  LAYER m7 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V7_120x40S_200H_120V

VIA V7_120x40S_200V_120V
  LAYER m7 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V7_120x40S_200V_120V

VIA V7_120x40S_80H_120V
  LAYER m7 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V7_120x40S_80H_120V

VIA V7_120x40_120H_120H
  LAYER m7 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V7_120x40_120H_120H

VIA V7_120x40_120H_160H
  LAYER m7 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V7_120x40_120H_160H

VIA V7_120x40_120H_160V
  LAYER m7 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V7_120x40_120H_160V

VIA V7_120x40_120H_200H
  LAYER m7 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V7_120x40_120H_200H

VIA V7_120x40_120H_200V
  LAYER m7 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V7_120x40_120H_200V

VIA V7_120x40_120H_80H
  LAYER m7 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V7_120x40_120H_80H

VIA V7_120x40_160H_120H
  LAYER m7 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V7_120x40_160H_120H

VIA V7_120x40_160H_160H
  LAYER m7 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V7_120x40_160H_160H

VIA V7_120x40_160H_160V
  LAYER m7 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V7_120x40_160H_160V

VIA V7_120x40_160H_200H
  LAYER m7 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V7_120x40_160H_200H

VIA V7_120x40_160H_200V
  LAYER m7 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V7_120x40_160H_200V

VIA V7_120x40_160H_80H
  LAYER m7 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V7_120x40_160H_80H

VIA V7_120x40_160V_120H
  LAYER m7 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V7_120x40_160V_120H

VIA V7_120x40_160V_160H
  LAYER m7 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V7_120x40_160V_160H

VIA V7_120x40_160V_160V
  LAYER m7 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V7_120x40_160V_160V

VIA V7_120x40_160V_200H
  LAYER m7 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V7_120x40_160V_200H

VIA V7_120x40_160V_200V
  LAYER m7 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V7_120x40_160V_200V

VIA V7_120x40_160V_80H
  LAYER m7 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V7_120x40_160V_80H

VIA V7_120x40_200H_120H
  LAYER m7 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V7_120x40_200H_120H

VIA V7_120x40_200H_160H
  LAYER m7 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V7_120x40_200H_160H

VIA V7_120x40_200H_160V
  LAYER m7 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V7_120x40_200H_160V

VIA V7_120x40_200H_200H
  LAYER m7 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V7_120x40_200H_200H

VIA V7_120x40_200H_200V
  LAYER m7 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V7_120x40_200H_200V

VIA V7_120x40_200H_80H
  LAYER m7 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V7_120x40_200H_80H

VIA V7_120x40_200V_120H
  LAYER m7 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V7_120x40_200V_120H

VIA V7_120x40_200V_160H
  LAYER m7 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V7_120x40_200V_160H

VIA V7_120x40_200V_160V
  LAYER m7 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V7_120x40_200V_160V

VIA V7_120x40_200V_200H
  LAYER m7 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V7_120x40_200V_200H

VIA V7_120x40_200V_200V
  LAYER m7 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V7_120x40_200V_200V

VIA V7_120x40_200V_80H
  LAYER m7 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V7_120x40_200V_80H

VIA V7_120x40_80H_120H
  LAYER m7 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V7_120x40_80H_120H

VIA V7_120x40_80H_160H
  LAYER m7 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V7_120x40_80H_160H

VIA V7_120x40_80H_160V
  LAYER m7 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V7_120x40_80H_160V

VIA V7_120x40_80H_200H
  LAYER m7 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V7_120x40_80H_200H

VIA V7_120x40_80H_200V
  LAYER m7 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V7_120x40_80H_200V

VIA V7_120x40_80H_80H
  LAYER m7 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v7 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m8 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V7_120x40_80H_80H

VIA V7_40Sx120_120H_120H
  LAYER m7 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V7_40Sx120_120H_120H

VIA V7_40Sx120_120V_120H
  LAYER m7 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V7_40Sx120_120V_120H

VIA V7_40Sx120_160H_120H
  LAYER m7 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V7_40Sx120_160H_120H

VIA V7_40Sx120_160V_120H
  LAYER m7 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V7_40Sx120_160V_120H

VIA V7_40Sx120_200H_120H
  LAYER m7 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V7_40Sx120_200H_120H

VIA V7_40Sx120_200V_120H
  LAYER m7 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V7_40Sx120_200V_120H

VIA V7_40Sx120_40V_120H
  LAYER m7 ;
    RECT -0.02 -0.084 0.02 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V7_40Sx120_40V_120H

VIA V7_40Sx120_60V_120H
  LAYER m7 ;
    RECT -0.03 -0.084 0.03 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V7_40Sx120_60V_120H

VIA V7_40Sx120_80V_120H
  LAYER m7 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V7_40Sx120_80V_120H

VIA V7_40Sx40_120H_40H
  LAYER m7 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v7 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m8 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V7_40Sx40_120H_40H

VIA V7_40Sx40_120V_40H
  LAYER m7 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v7 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m8 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V7_40Sx40_120V_40H

VIA V7_40Sx40_160H_40H
  LAYER m7 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v7 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m8 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V7_40Sx40_160H_40H

VIA V7_40Sx40_160V_40H
  LAYER m7 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v7 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m8 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V7_40Sx40_160V_40H

VIA V7_40Sx40_200H_40H
  LAYER m7 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v7 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m8 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V7_40Sx40_200H_40H

VIA V7_40Sx40_200V_40H
  LAYER m7 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v7 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m8 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V7_40Sx40_200V_40H

VIA V7_40Sx40_40V_40H
  LAYER m7 ;
    RECT -0.02 -0.044 0.02 0.044 ;
  LAYER v7 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m8 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V7_40Sx40_40V_40H

VIA V7_40Sx40_60V_40H
  LAYER m7 ;
    RECT -0.03 -0.044 0.03 0.044 ;
  LAYER v7 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m8 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V7_40Sx40_60V_40H

VIA V7_40Sx40_80H_40H
  LAYER m7 ;
    RECT -0.044 -0.04 0.044 0.04 ;
  LAYER v7 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m8 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V7_40Sx40_80H_40H

VIA V7_40Sx40_80V_40H
  LAYER m7 ;
    RECT -0.04 -0.044 0.04 0.044 ;
  LAYER v7 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m8 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V7_40Sx40_80V_40H

VIA V7_40Sx60_120H_60H
  LAYER m7 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v7 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m8 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V7_40Sx60_120H_60H

VIA V7_40Sx60_120V_60H
  LAYER m7 ;
    RECT -0.06 -0.054 0.06 0.054 ;
  LAYER v7 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m8 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V7_40Sx60_120V_60H

VIA V7_40Sx60_160H_60H
  LAYER m7 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v7 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m8 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V7_40Sx60_160H_60H

VIA V7_40Sx60_160V_60H
  LAYER m7 ;
    RECT -0.08 -0.054 0.08 0.054 ;
  LAYER v7 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m8 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V7_40Sx60_160V_60H

VIA V7_40Sx60_200H_60H
  LAYER m7 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v7 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m8 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V7_40Sx60_200H_60H

VIA V7_40Sx60_200V_60H
  LAYER m7 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v7 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m8 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V7_40Sx60_200V_60H

VIA V7_40Sx60_40V_60H
  LAYER m7 ;
    RECT -0.02 -0.054 0.02 0.054 ;
  LAYER v7 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m8 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V7_40Sx60_40V_60H

VIA V7_40Sx60_60V_60H
  LAYER m7 ;
    RECT -0.03 -0.054 0.03 0.054 ;
  LAYER v7 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m8 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V7_40Sx60_60V_60H

VIA V7_40Sx60_80H_60H
  LAYER m7 ;
    RECT -0.044 -0.04 0.044 0.04 ;
  LAYER v7 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m8 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V7_40Sx60_80H_60H

VIA V7_40Sx60_80V_60H
  LAYER m7 ;
    RECT -0.04 -0.054 0.04 0.054 ;
  LAYER v7 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m8 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V7_40Sx60_80V_60H

VIA V7_40Sx80_120H_80H
  LAYER m7 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v7 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m8 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V7_40Sx80_120H_80H

VIA V7_40Sx80_120V_80H
  LAYER m7 ;
    RECT -0.06 -0.064 0.06 0.064 ;
  LAYER v7 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m8 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V7_40Sx80_120V_80H

VIA V7_40Sx80_160H_80H
  LAYER m7 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v7 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m8 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V7_40Sx80_160H_80H

VIA V7_40Sx80_160V_80H
  LAYER m7 ;
    RECT -0.08 -0.064 0.08 0.064 ;
  LAYER v7 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m8 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V7_40Sx80_160V_80H

VIA V7_40Sx80_200H_80H
  LAYER m7 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v7 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m8 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V7_40Sx80_200H_80H

VIA V7_40Sx80_200V_80H
  LAYER m7 ;
    RECT -0.1 -0.064 0.1 0.064 ;
  LAYER v7 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m8 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V7_40Sx80_200V_80H

VIA V7_40Sx80_40V_80H
  LAYER m7 ;
    RECT -0.02 -0.064 0.02 0.064 ;
  LAYER v7 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m8 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V7_40Sx80_40V_80H

VIA V7_40Sx80_60V_80H
  LAYER m7 ;
    RECT -0.03 -0.064 0.03 0.064 ;
  LAYER v7 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m8 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V7_40Sx80_60V_80H

VIA V7_40Sx80_80H_80H
  LAYER m7 ;
    RECT -0.044 -0.04 0.044 0.04 ;
  LAYER v7 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m8 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V7_40Sx80_80H_80H

VIA V7_40Sx80_80V_80H
  LAYER m7 ;
    RECT -0.04 -0.064 0.04 0.064 ;
  LAYER v7 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m8 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V7_40Sx80_80V_80H

VIA V7_40x120_120V_120V
  LAYER m7 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V7_40x120_120V_120V

VIA V7_40x120_120V_160H
  LAYER m7 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V7_40x120_120V_160H

VIA V7_40x120_120V_160V
  LAYER m7 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V7_40x120_120V_160V

VIA V7_40x120_120V_200H
  LAYER m7 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V7_40x120_120V_200H

VIA V7_40x120_120V_200V
  LAYER m7 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V7_40x120_120V_200V

VIA V7_40x120_120V_80V
  LAYER m7 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V7_40x120_120V_80V

VIA V7_40x120_160H_120V
  LAYER m7 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V7_40x120_160H_120V

VIA V7_40x120_160H_160H
  LAYER m7 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V7_40x120_160H_160H

VIA V7_40x120_160H_160V
  LAYER m7 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V7_40x120_160H_160V

VIA V7_40x120_160H_200H
  LAYER m7 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V7_40x120_160H_200H

VIA V7_40x120_160H_200V
  LAYER m7 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V7_40x120_160H_200V

VIA V7_40x120_160H_80V
  LAYER m7 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V7_40x120_160H_80V

VIA V7_40x120_160V_120V
  LAYER m7 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V7_40x120_160V_120V

VIA V7_40x120_160V_160H
  LAYER m7 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V7_40x120_160V_160H

VIA V7_40x120_160V_160V
  LAYER m7 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V7_40x120_160V_160V

VIA V7_40x120_160V_200H
  LAYER m7 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V7_40x120_160V_200H

VIA V7_40x120_160V_200V
  LAYER m7 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V7_40x120_160V_200V

VIA V7_40x120_160V_80V
  LAYER m7 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V7_40x120_160V_80V

VIA V7_40x120_200H_120V
  LAYER m7 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V7_40x120_200H_120V

VIA V7_40x120_200H_160H
  LAYER m7 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V7_40x120_200H_160H

VIA V7_40x120_200H_160V
  LAYER m7 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V7_40x120_200H_160V

VIA V7_40x120_200H_200H
  LAYER m7 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V7_40x120_200H_200H

VIA V7_40x120_200H_200V
  LAYER m7 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V7_40x120_200H_200V

VIA V7_40x120_200H_80V
  LAYER m7 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V7_40x120_200H_80V

VIA V7_40x120_200V_120V
  LAYER m7 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V7_40x120_200V_120V

VIA V7_40x120_200V_160H
  LAYER m7 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V7_40x120_200V_160H

VIA V7_40x120_200V_160V
  LAYER m7 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V7_40x120_200V_160V

VIA V7_40x120_200V_200H
  LAYER m7 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V7_40x120_200V_200H

VIA V7_40x120_200V_200V
  LAYER m7 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V7_40x120_200V_200V

VIA V7_40x120_200V_80V
  LAYER m7 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V7_40x120_200V_80V

VIA V7_40x120_80V_120V
  LAYER m7 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V7_40x120_80V_120V

VIA V7_40x120_80V_160H
  LAYER m7 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V7_40x120_80V_160H

VIA V7_40x120_80V_160V
  LAYER m7 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V7_40x120_80V_160V

VIA V7_40x120_80V_200H
  LAYER m7 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V7_40x120_80V_200H

VIA V7_40x120_80V_200V
  LAYER m7 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V7_40x120_80V_200V

VIA V7_40x120_80V_80V
  LAYER m7 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v7 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m8 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V7_40x120_80V_80V

VIA V7_60Sx40_120H_40H
  LAYER m7 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v7 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m8 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V7_60Sx40_120H_40H

VIA V7_60Sx40_120V_40H
  LAYER m7 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v7 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m8 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V7_60Sx40_120V_40H

VIA V7_60Sx40_160H_40H
  LAYER m7 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v7 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m8 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V7_60Sx40_160H_40H

VIA V7_60Sx40_160V_40H
  LAYER m7 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v7 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m8 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V7_60Sx40_160V_40H

VIA V7_60Sx40_200H_40H
  LAYER m7 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v7 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m8 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V7_60Sx40_200H_40H

VIA V7_60Sx40_200V_40H
  LAYER m7 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v7 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m8 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V7_60Sx40_200V_40H

VIA V7_60Sx40_60V_40H
  LAYER m7 ;
    RECT -0.03 -0.044 0.03 0.044 ;
  LAYER v7 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m8 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V7_60Sx40_60V_40H

VIA V7_60Sx40_80H_40H
  LAYER m7 ;
    RECT -0.054 -0.04 0.054 0.04 ;
  LAYER v7 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m8 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V7_60Sx40_80H_40H

VIA V7_60Sx40_80V_40H
  LAYER m7 ;
    RECT -0.04 -0.044 0.04 0.044 ;
  LAYER v7 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m8 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V7_60Sx40_80V_40H

VIA V7_60Sx60_120H_60H
  LAYER m7 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v7 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m8 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V7_60Sx60_120H_60H

VIA V7_60Sx60_120V_60H
  LAYER m7 ;
    RECT -0.06 -0.054 0.06 0.054 ;
  LAYER v7 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m8 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V7_60Sx60_120V_60H

VIA V7_60Sx60_160H_60H
  LAYER m7 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v7 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m8 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V7_60Sx60_160H_60H

VIA V7_60Sx60_160V_60H
  LAYER m7 ;
    RECT -0.08 -0.054 0.08 0.054 ;
  LAYER v7 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m8 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V7_60Sx60_160V_60H

VIA V7_60Sx60_200H_60H
  LAYER m7 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v7 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m8 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V7_60Sx60_200H_60H

VIA V7_60Sx60_200V_60H
  LAYER m7 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v7 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m8 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V7_60Sx60_200V_60H

VIA V7_60Sx60_60V_60H
  LAYER m7 ;
    RECT -0.03 -0.054 0.03 0.054 ;
  LAYER v7 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m8 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V7_60Sx60_60V_60H

VIA V7_60Sx60_80H_60H
  LAYER m7 ;
    RECT -0.054 -0.04 0.054 0.04 ;
  LAYER v7 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m8 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V7_60Sx60_80H_60H

VIA V7_60Sx60_80V_60H
  LAYER m7 ;
    RECT -0.04 -0.054 0.04 0.054 ;
  LAYER v7 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m8 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V7_60Sx60_80V_60H

VIA V7_60Sx80_120H_80H
  LAYER m7 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v7 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m8 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V7_60Sx80_120H_80H

VIA V7_60Sx80_120V_80H
  LAYER m7 ;
    RECT -0.06 -0.064 0.06 0.064 ;
  LAYER v7 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m8 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V7_60Sx80_120V_80H

VIA V7_60Sx80_160H_80H
  LAYER m7 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v7 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m8 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V7_60Sx80_160H_80H

VIA V7_60Sx80_160V_80H
  LAYER m7 ;
    RECT -0.08 -0.064 0.08 0.064 ;
  LAYER v7 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m8 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V7_60Sx80_160V_80H

VIA V7_60Sx80_200H_80H
  LAYER m7 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v7 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m8 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V7_60Sx80_200H_80H

VIA V7_60Sx80_200V_80H
  LAYER m7 ;
    RECT -0.1 -0.064 0.1 0.064 ;
  LAYER v7 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m8 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V7_60Sx80_200V_80H

VIA V7_60Sx80_60V_80H
  LAYER m7 ;
    RECT -0.03 -0.064 0.03 0.064 ;
  LAYER v7 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m8 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V7_60Sx80_60V_80H

VIA V7_60Sx80_80H_80H
  LAYER m7 ;
    RECT -0.054 -0.04 0.054 0.04 ;
  LAYER v7 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m8 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V7_60Sx80_80H_80H

VIA V7_60Sx80_80V_80H
  LAYER m7 ;
    RECT -0.04 -0.064 0.04 0.064 ;
  LAYER v7 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m8 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V7_60Sx80_80V_80H

VIA V7_80x40S_120H_80V
  LAYER m7 ;
    RECT -0.064 -0.06 0.064 0.06 ;
  LAYER v7 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m8 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V7_80x40S_120H_80V

VIA V7_80x40S_120V_80V
  LAYER m7 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v7 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m8 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V7_80x40S_120V_80V

VIA V7_80x40S_160H_80V
  LAYER m7 ;
    RECT -0.064 -0.08 0.064 0.08 ;
  LAYER v7 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m8 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V7_80x40S_160H_80V

VIA V7_80x40S_160V_80V
  LAYER m7 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v7 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m8 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V7_80x40S_160V_80V

VIA V7_80x40S_200H_80V
  LAYER m7 ;
    RECT -0.064 -0.1 0.064 0.1 ;
  LAYER v7 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m8 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V7_80x40S_200H_80V

VIA V7_80x40S_200V_80V
  LAYER m7 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v7 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m8 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V7_80x40S_200V_80V

VIA V7_80x40S_80H_80V
  LAYER m7 ;
    RECT -0.064 -0.04 0.064 0.04 ;
  LAYER v7 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m8 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V7_80x40S_80H_80V

VIA V7_80x40S_80V_80V
  LAYER m7 ;
    RECT -0.04 -0.044 0.04 0.044 ;
  LAYER v7 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m8 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V7_80x40S_80V_80V

VIA V8_120x40S_120H_120V
  LAYER m8 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V8_120x40S_120H_120V

VIA V8_120x40S_120V_120V
  LAYER m8 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V8_120x40S_120V_120V

VIA V8_120x40S_160H_120V
  LAYER m8 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V8_120x40S_160H_120V

VIA V8_120x40S_160V_120V
  LAYER m8 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V8_120x40S_160V_120V

VIA V8_120x40S_200H_120V
  LAYER m8 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V8_120x40S_200H_120V

VIA V8_120x40S_200V_120V
  LAYER m8 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V8_120x40S_200V_120V

VIA V8_120x40S_40H_120V
  LAYER m8 ;
    RECT -0.084 -0.02 0.084 0.02 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V8_120x40S_40H_120V

VIA V8_120x40S_60H_120V
  LAYER m8 ;
    RECT -0.084 -0.03 0.084 0.03 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V8_120x40S_60H_120V

VIA V8_120x40S_80H_120V
  LAYER m8 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V8_120x40S_80H_120V

VIA V8_120x40_120H_120H
  LAYER m8 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V8_120x40_120H_120H

VIA V8_120x40_120H_160H
  LAYER m8 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V8_120x40_120H_160H

VIA V8_120x40_120H_160V
  LAYER m8 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V8_120x40_120H_160V

VIA V8_120x40_120H_200H
  LAYER m8 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V8_120x40_120H_200H

VIA V8_120x40_120H_200V
  LAYER m8 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V8_120x40_120H_200V

VIA V8_120x40_120H_80H
  LAYER m8 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V8_120x40_120H_80H

VIA V8_120x40_160H_120H
  LAYER m8 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V8_120x40_160H_120H

VIA V8_120x40_160H_160H
  LAYER m8 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V8_120x40_160H_160H

VIA V8_120x40_160H_160V
  LAYER m8 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V8_120x40_160H_160V

VIA V8_120x40_160H_200H
  LAYER m8 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V8_120x40_160H_200H

VIA V8_120x40_160H_200V
  LAYER m8 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V8_120x40_160H_200V

VIA V8_120x40_160H_80H
  LAYER m8 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V8_120x40_160H_80H

VIA V8_120x40_160V_120H
  LAYER m8 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V8_120x40_160V_120H

VIA V8_120x40_160V_160H
  LAYER m8 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V8_120x40_160V_160H

VIA V8_120x40_160V_160V
  LAYER m8 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V8_120x40_160V_160V

VIA V8_120x40_160V_200H
  LAYER m8 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V8_120x40_160V_200H

VIA V8_120x40_160V_200V
  LAYER m8 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V8_120x40_160V_200V

VIA V8_120x40_160V_80H
  LAYER m8 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V8_120x40_160V_80H

VIA V8_120x40_200H_120H
  LAYER m8 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V8_120x40_200H_120H

VIA V8_120x40_200H_160H
  LAYER m8 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V8_120x40_200H_160H

VIA V8_120x40_200H_160V
  LAYER m8 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V8_120x40_200H_160V

VIA V8_120x40_200H_200H
  LAYER m8 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V8_120x40_200H_200H

VIA V8_120x40_200H_200V
  LAYER m8 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V8_120x40_200H_200V

VIA V8_120x40_200H_80H
  LAYER m8 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V8_120x40_200H_80H

VIA V8_120x40_200V_120H
  LAYER m8 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V8_120x40_200V_120H

VIA V8_120x40_200V_160H
  LAYER m8 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V8_120x40_200V_160H

VIA V8_120x40_200V_160V
  LAYER m8 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V8_120x40_200V_160V

VIA V8_120x40_200V_200H
  LAYER m8 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V8_120x40_200V_200H

VIA V8_120x40_200V_200V
  LAYER m8 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V8_120x40_200V_200V

VIA V8_120x40_200V_80H
  LAYER m8 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V8_120x40_200V_80H

VIA V8_120x40_80H_120H
  LAYER m8 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V8_120x40_80H_120H

VIA V8_120x40_80H_160H
  LAYER m8 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V8_120x40_80H_160H

VIA V8_120x40_80H_160V
  LAYER m8 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V8_120x40_80H_160V

VIA V8_120x40_80H_200H
  LAYER m8 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V8_120x40_80H_200H

VIA V8_120x40_80H_200V
  LAYER m8 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V8_120x40_80H_200V

VIA V8_120x40_80H_80H
  LAYER m8 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v8 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m9 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V8_120x40_80H_80H

VIA V8_40Sx120_120H_120H
  LAYER m8 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V8_40Sx120_120H_120H

VIA V8_40Sx120_120V_120H
  LAYER m8 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V8_40Sx120_120V_120H

VIA V8_40Sx120_160H_120H
  LAYER m8 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V8_40Sx120_160H_120H

VIA V8_40Sx120_160V_120H
  LAYER m8 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V8_40Sx120_160V_120H

VIA V8_40Sx120_200H_120H
  LAYER m8 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V8_40Sx120_200H_120H

VIA V8_40Sx120_200V_120H
  LAYER m8 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V8_40Sx120_200V_120H

VIA V8_40Sx120_80V_120H
  LAYER m8 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V8_40Sx120_80V_120H

VIA V8_40Sx80_120H_80H
  LAYER m8 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v8 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m9 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V8_40Sx80_120H_80H

VIA V8_40Sx80_120V_80H
  LAYER m8 ;
    RECT -0.06 -0.064 0.06 0.064 ;
  LAYER v8 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m9 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V8_40Sx80_120V_80H

VIA V8_40Sx80_160H_80H
  LAYER m8 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v8 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m9 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V8_40Sx80_160H_80H

VIA V8_40Sx80_160V_80H
  LAYER m8 ;
    RECT -0.08 -0.064 0.08 0.064 ;
  LAYER v8 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m9 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V8_40Sx80_160V_80H

VIA V8_40Sx80_200H_80H
  LAYER m8 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v8 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m9 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V8_40Sx80_200H_80H

VIA V8_40Sx80_200V_80H
  LAYER m8 ;
    RECT -0.1 -0.064 0.1 0.064 ;
  LAYER v8 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m9 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V8_40Sx80_200V_80H

VIA V8_40Sx80_80H_80H
  LAYER m8 ;
    RECT -0.044 -0.04 0.044 0.04 ;
  LAYER v8 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m9 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V8_40Sx80_80H_80H

VIA V8_40Sx80_80V_80H
  LAYER m8 ;
    RECT -0.04 -0.064 0.04 0.064 ;
  LAYER v8 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m9 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V8_40Sx80_80V_80H

VIA V8_40x120_120V_120V
  LAYER m8 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V8_40x120_120V_120V

VIA V8_40x120_120V_160H
  LAYER m8 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V8_40x120_120V_160H

VIA V8_40x120_120V_160V
  LAYER m8 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V8_40x120_120V_160V

VIA V8_40x120_120V_200H
  LAYER m8 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V8_40x120_120V_200H

VIA V8_40x120_120V_200V
  LAYER m8 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V8_40x120_120V_200V

VIA V8_40x120_120V_80V
  LAYER m8 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V8_40x120_120V_80V

VIA V8_40x120_160H_120V
  LAYER m8 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V8_40x120_160H_120V

VIA V8_40x120_160H_160H
  LAYER m8 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V8_40x120_160H_160H

VIA V8_40x120_160H_160V
  LAYER m8 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V8_40x120_160H_160V

VIA V8_40x120_160H_200H
  LAYER m8 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V8_40x120_160H_200H

VIA V8_40x120_160H_200V
  LAYER m8 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V8_40x120_160H_200V

VIA V8_40x120_160H_80V
  LAYER m8 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V8_40x120_160H_80V

VIA V8_40x120_160V_120V
  LAYER m8 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V8_40x120_160V_120V

VIA V8_40x120_160V_160H
  LAYER m8 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V8_40x120_160V_160H

VIA V8_40x120_160V_160V
  LAYER m8 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V8_40x120_160V_160V

VIA V8_40x120_160V_200H
  LAYER m8 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V8_40x120_160V_200H

VIA V8_40x120_160V_200V
  LAYER m8 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V8_40x120_160V_200V

VIA V8_40x120_160V_80V
  LAYER m8 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V8_40x120_160V_80V

VIA V8_40x120_200H_120V
  LAYER m8 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V8_40x120_200H_120V

VIA V8_40x120_200H_160H
  LAYER m8 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V8_40x120_200H_160H

VIA V8_40x120_200H_160V
  LAYER m8 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V8_40x120_200H_160V

VIA V8_40x120_200H_200H
  LAYER m8 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V8_40x120_200H_200H

VIA V8_40x120_200H_200V
  LAYER m8 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V8_40x120_200H_200V

VIA V8_40x120_200H_80V
  LAYER m8 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V8_40x120_200H_80V

VIA V8_40x120_200V_120V
  LAYER m8 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V8_40x120_200V_120V

VIA V8_40x120_200V_160H
  LAYER m8 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V8_40x120_200V_160H

VIA V8_40x120_200V_160V
  LAYER m8 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V8_40x120_200V_160V

VIA V8_40x120_200V_200H
  LAYER m8 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V8_40x120_200V_200H

VIA V8_40x120_200V_200V
  LAYER m8 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V8_40x120_200V_200V

VIA V8_40x120_200V_80V
  LAYER m8 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V8_40x120_200V_80V

VIA V8_40x120_80V_120V
  LAYER m8 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V8_40x120_80V_120V

VIA V8_40x120_80V_160H
  LAYER m8 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V8_40x120_80V_160H

VIA V8_40x120_80V_160V
  LAYER m8 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V8_40x120_80V_160V

VIA V8_40x120_80V_200H
  LAYER m8 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V8_40x120_80V_200H

VIA V8_40x120_80V_200V
  LAYER m8 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V8_40x120_80V_200V

VIA V8_40x120_80V_80V
  LAYER m8 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v8 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m9 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V8_40x120_80V_80V

VIA V8_40x40S_120H_40V
  LAYER m8 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v8 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m9 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V8_40x40S_120H_40V

VIA V8_40x40S_120V_40V
  LAYER m8 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v8 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m9 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V8_40x40S_120V_40V

VIA V8_40x40S_160H_40V
  LAYER m8 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v8 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m9 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V8_40x40S_160H_40V

VIA V8_40x40S_160V_40V
  LAYER m8 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v8 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m9 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V8_40x40S_160V_40V

VIA V8_40x40S_200H_40V
  LAYER m8 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v8 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m9 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V8_40x40S_200H_40V

VIA V8_40x40S_200V_40V
  LAYER m8 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v8 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m9 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V8_40x40S_200V_40V

VIA V8_40x40S_40H_40V
  LAYER m8 ;
    RECT -0.044 -0.02 0.044 0.02 ;
  LAYER v8 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m9 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V8_40x40S_40H_40V

VIA V8_40x40S_60H_40V
  LAYER m8 ;
    RECT -0.044 -0.03 0.044 0.03 ;
  LAYER v8 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m9 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V8_40x40S_60H_40V

VIA V8_40x40S_80H_40V
  LAYER m8 ;
    RECT -0.044 -0.04 0.044 0.04 ;
  LAYER v8 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m9 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V8_40x40S_80H_40V

VIA V8_40x40S_80V_40V
  LAYER m8 ;
    RECT -0.04 -0.044 0.04 0.044 ;
  LAYER v8 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m9 ;
    RECT -0.02 -0.058 0.02 0.058 ;
END V8_40x40S_80V_40V

VIA V8_40x60S_120H_40V
  LAYER m8 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v8 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m9 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V8_40x60S_120H_40V

VIA V8_40x60S_120V_40V
  LAYER m8 ;
    RECT -0.06 -0.054 0.06 0.054 ;
  LAYER v8 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m9 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V8_40x60S_120V_40V

VIA V8_40x60S_160H_40V
  LAYER m8 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v8 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m9 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V8_40x60S_160H_40V

VIA V8_40x60S_160V_40V
  LAYER m8 ;
    RECT -0.08 -0.054 0.08 0.054 ;
  LAYER v8 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m9 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V8_40x60S_160V_40V

VIA V8_40x60S_200H_40V
  LAYER m8 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v8 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m9 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V8_40x60S_200H_40V

VIA V8_40x60S_200V_40V
  LAYER m8 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v8 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m9 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V8_40x60S_200V_40V

VIA V8_40x60S_60H_40V
  LAYER m8 ;
    RECT -0.044 -0.03 0.044 0.03 ;
  LAYER v8 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m9 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V8_40x60S_60H_40V

VIA V8_40x60S_80H_40V
  LAYER m8 ;
    RECT -0.044 -0.04 0.044 0.04 ;
  LAYER v8 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m9 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V8_40x60S_80H_40V

VIA V8_40x60S_80V_40V
  LAYER m8 ;
    RECT -0.04 -0.054 0.04 0.054 ;
  LAYER v8 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m9 ;
    RECT -0.02 -0.068 0.02 0.068 ;
END V8_40x60S_80V_40V

VIA V8_60x40S_120H_60V
  LAYER m8 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v8 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m9 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V8_60x40S_120H_60V

VIA V8_60x40S_120V_60V
  LAYER m8 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v8 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m9 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V8_60x40S_120V_60V

VIA V8_60x40S_160H_60V
  LAYER m8 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v8 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m9 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V8_60x40S_160H_60V

VIA V8_60x40S_160V_60V
  LAYER m8 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v8 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m9 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V8_60x40S_160V_60V

VIA V8_60x40S_200H_60V
  LAYER m8 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v8 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m9 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V8_60x40S_200H_60V

VIA V8_60x40S_200V_60V
  LAYER m8 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v8 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m9 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V8_60x40S_200V_60V

VIA V8_60x40S_40H_60V
  LAYER m8 ;
    RECT -0.054 -0.02 0.054 0.02 ;
  LAYER v8 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m9 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V8_60x40S_40H_60V

VIA V8_60x40S_60H_60V
  LAYER m8 ;
    RECT -0.054 -0.03 0.054 0.03 ;
  LAYER v8 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m9 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V8_60x40S_60H_60V

VIA V8_60x40S_80H_60V
  LAYER m8 ;
    RECT -0.054 -0.04 0.054 0.04 ;
  LAYER v8 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m9 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V8_60x40S_80H_60V

VIA V8_60x40S_80V_60V
  LAYER m8 ;
    RECT -0.04 -0.044 0.04 0.044 ;
  LAYER v8 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m9 ;
    RECT -0.03 -0.058 0.03 0.058 ;
END V8_60x40S_80V_60V

VIA V8_60x60S_120H_60V
  LAYER m8 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v8 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m9 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V8_60x60S_120H_60V

VIA V8_60x60S_120V_60V
  LAYER m8 ;
    RECT -0.06 -0.054 0.06 0.054 ;
  LAYER v8 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m9 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V8_60x60S_120V_60V

VIA V8_60x60S_160H_60V
  LAYER m8 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v8 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m9 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V8_60x60S_160H_60V

VIA V8_60x60S_160V_60V
  LAYER m8 ;
    RECT -0.08 -0.054 0.08 0.054 ;
  LAYER v8 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m9 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V8_60x60S_160V_60V

VIA V8_60x60S_200H_60V
  LAYER m8 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v8 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m9 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V8_60x60S_200H_60V

VIA V8_60x60S_200V_60V
  LAYER m8 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v8 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m9 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V8_60x60S_200V_60V

VIA V8_60x60S_60H_60V
  LAYER m8 ;
    RECT -0.054 -0.03 0.054 0.03 ;
  LAYER v8 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m9 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V8_60x60S_60H_60V

VIA V8_60x60S_80H_60V
  LAYER m8 ;
    RECT -0.054 -0.04 0.054 0.04 ;
  LAYER v8 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m9 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V8_60x60S_80H_60V

VIA V8_60x60S_80V_60V
  LAYER m8 ;
    RECT -0.04 -0.054 0.04 0.054 ;
  LAYER v8 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m9 ;
    RECT -0.03 -0.068 0.03 0.068 ;
END V8_60x60S_80V_60V

VIA V8_80x40S_120H_80V
  LAYER m8 ;
    RECT -0.064 -0.06 0.064 0.06 ;
  LAYER v8 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m9 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V8_80x40S_120H_80V

VIA V8_80x40S_120V_80V
  LAYER m8 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v8 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m9 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V8_80x40S_120V_80V

VIA V8_80x40S_160H_80V
  LAYER m8 ;
    RECT -0.064 -0.08 0.064 0.08 ;
  LAYER v8 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m9 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V8_80x40S_160H_80V

VIA V8_80x40S_160V_80V
  LAYER m8 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v8 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m9 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V8_80x40S_160V_80V

VIA V8_80x40S_200H_80V
  LAYER m8 ;
    RECT -0.064 -0.1 0.064 0.1 ;
  LAYER v8 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m9 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V8_80x40S_200H_80V

VIA V8_80x40S_200V_80V
  LAYER m8 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v8 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m9 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V8_80x40S_200V_80V

VIA V8_80x40S_40H_80V
  LAYER m8 ;
    RECT -0.064 -0.02 0.064 0.02 ;
  LAYER v8 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m9 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V8_80x40S_40H_80V

VIA V8_80x40S_60H_80V
  LAYER m8 ;
    RECT -0.064 -0.03 0.064 0.03 ;
  LAYER v8 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m9 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V8_80x40S_60H_80V

VIA V8_80x40S_80H_80V
  LAYER m8 ;
    RECT -0.064 -0.04 0.064 0.04 ;
  LAYER v8 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m9 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V8_80x40S_80H_80V

VIA V8_80x40S_80V_80V
  LAYER m8 ;
    RECT -0.04 -0.044 0.04 0.044 ;
  LAYER v8 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m9 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V8_80x40S_80V_80V

VIA V8_80x60S_120H_80V
  LAYER m8 ;
    RECT -0.064 -0.06 0.064 0.06 ;
  LAYER v8 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m9 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V8_80x60S_120H_80V

VIA V8_80x60S_120V_80V
  LAYER m8 ;
    RECT -0.06 -0.054 0.06 0.054 ;
  LAYER v8 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m9 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V8_80x60S_120V_80V

VIA V8_80x60S_160H_80V
  LAYER m8 ;
    RECT -0.064 -0.08 0.064 0.08 ;
  LAYER v8 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m9 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V8_80x60S_160H_80V

VIA V8_80x60S_160V_80V
  LAYER m8 ;
    RECT -0.08 -0.054 0.08 0.054 ;
  LAYER v8 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m9 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V8_80x60S_160V_80V

VIA V8_80x60S_200H_80V
  LAYER m8 ;
    RECT -0.064 -0.1 0.064 0.1 ;
  LAYER v8 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m9 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V8_80x60S_200H_80V

VIA V8_80x60S_200V_80V
  LAYER m8 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v8 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m9 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V8_80x60S_200V_80V

VIA V8_80x60S_60H_80V
  LAYER m8 ;
    RECT -0.064 -0.03 0.064 0.03 ;
  LAYER v8 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m9 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V8_80x60S_60H_80V

VIA V8_80x60S_80H_80V
  LAYER m8 ;
    RECT -0.064 -0.04 0.064 0.04 ;
  LAYER v8 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m9 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V8_80x60S_80H_80V

VIA V8_80x60S_80V_80V
  LAYER m8 ;
    RECT -0.04 -0.054 0.04 0.054 ;
  LAYER v8 ;
    RECT -0.04 -0.03 0.04 0.03 ;
  LAYER m9 ;
    RECT -0.04 -0.068 0.04 0.068 ;
END V8_80x60S_80V_80V

VIA V9_120x40S_120H_120V
  LAYER m9 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V9_120x40S_120H_120V

VIA V9_120x40S_120V_120V
  LAYER m9 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V9_120x40S_120V_120V

VIA V9_120x40S_160H_120V
  LAYER m9 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V9_120x40S_160H_120V

VIA V9_120x40S_160V_120V
  LAYER m9 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V9_120x40S_160V_120V

VIA V9_120x40S_200H_120V
  LAYER m9 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V9_120x40S_200H_120V

VIA V9_120x40S_200V_120V
  LAYER m9 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V9_120x40S_200V_120V

VIA V9_120x40S_80H_120V
  LAYER m9 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.06 -0.058 0.06 0.058 ;
END V9_120x40S_80H_120V

VIA V9_120x40_120H_120H
  LAYER m9 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V9_120x40_120H_120H

VIA V9_120x40_120H_160H
  LAYER m9 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V9_120x40_120H_160H

VIA V9_120x40_120H_160V
  LAYER m9 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V9_120x40_120H_160V

VIA V9_120x40_120H_200H
  LAYER m9 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V9_120x40_120H_200H

VIA V9_120x40_120H_200V
  LAYER m9 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V9_120x40_120H_200V

VIA V9_120x40_120H_80H
  LAYER m9 ;
    RECT -0.084 -0.06 0.084 0.06 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V9_120x40_120H_80H

VIA V9_120x40_160H_120H
  LAYER m9 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V9_120x40_160H_120H

VIA V9_120x40_160H_160H
  LAYER m9 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V9_120x40_160H_160H

VIA V9_120x40_160H_160V
  LAYER m9 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V9_120x40_160H_160V

VIA V9_120x40_160H_200H
  LAYER m9 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V9_120x40_160H_200H

VIA V9_120x40_160H_200V
  LAYER m9 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V9_120x40_160H_200V

VIA V9_120x40_160H_80H
  LAYER m9 ;
    RECT -0.084 -0.08 0.084 0.08 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V9_120x40_160H_80H

VIA V9_120x40_160V_120H
  LAYER m9 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V9_120x40_160V_120H

VIA V9_120x40_160V_160H
  LAYER m9 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V9_120x40_160V_160H

VIA V9_120x40_160V_160V
  LAYER m9 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V9_120x40_160V_160V

VIA V9_120x40_160V_200H
  LAYER m9 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V9_120x40_160V_200H

VIA V9_120x40_160V_200V
  LAYER m9 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V9_120x40_160V_200V

VIA V9_120x40_160V_80H
  LAYER m9 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V9_120x40_160V_80H

VIA V9_120x40_200H_120H
  LAYER m9 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V9_120x40_200H_120H

VIA V9_120x40_200H_160H
  LAYER m9 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V9_120x40_200H_160H

VIA V9_120x40_200H_160V
  LAYER m9 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V9_120x40_200H_160V

VIA V9_120x40_200H_200H
  LAYER m9 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V9_120x40_200H_200H

VIA V9_120x40_200H_200V
  LAYER m9 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V9_120x40_200H_200V

VIA V9_120x40_200H_80H
  LAYER m9 ;
    RECT -0.084 -0.1 0.084 0.1 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V9_120x40_200H_80H

VIA V9_120x40_200V_120H
  LAYER m9 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V9_120x40_200V_120H

VIA V9_120x40_200V_160H
  LAYER m9 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V9_120x40_200V_160H

VIA V9_120x40_200V_160V
  LAYER m9 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V9_120x40_200V_160V

VIA V9_120x40_200V_200H
  LAYER m9 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V9_120x40_200V_200H

VIA V9_120x40_200V_200V
  LAYER m9 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V9_120x40_200V_200V

VIA V9_120x40_200V_80H
  LAYER m9 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V9_120x40_200V_80H

VIA V9_120x40_80H_120H
  LAYER m9 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.06 0.098 0.06 ;
END V9_120x40_80H_120H

VIA V9_120x40_80H_160H
  LAYER m9 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.08 0.098 0.08 ;
END V9_120x40_80H_160H

VIA V9_120x40_80H_160V
  LAYER m9 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.08 -0.058 0.08 0.058 ;
END V9_120x40_80H_160V

VIA V9_120x40_80H_200H
  LAYER m9 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.1 0.098 0.1 ;
END V9_120x40_80H_200H

VIA V9_120x40_80H_200V
  LAYER m9 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.1 -0.058 0.1 0.058 ;
END V9_120x40_80H_200V

VIA V9_120x40_80H_80H
  LAYER m9 ;
    RECT -0.084 -0.04 0.084 0.04 ;
  LAYER v9 ;
    RECT -0.06 -0.02 0.06 0.02 ;
  LAYER m10 ;
    RECT -0.098 -0.04 0.098 0.04 ;
END V9_120x40_80H_80H

VIA V9_40Sx120_120H_120H
  LAYER m9 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V9_40Sx120_120H_120H

VIA V9_40Sx120_120V_120H
  LAYER m9 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V9_40Sx120_120V_120H

VIA V9_40Sx120_160H_120H
  LAYER m9 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V9_40Sx120_160H_120H

VIA V9_40Sx120_160V_120H
  LAYER m9 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V9_40Sx120_160V_120H

VIA V9_40Sx120_200H_120H
  LAYER m9 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V9_40Sx120_200H_120H

VIA V9_40Sx120_200V_120H
  LAYER m9 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V9_40Sx120_200V_120H

VIA V9_40Sx120_40V_120H
  LAYER m9 ;
    RECT -0.02 -0.084 0.02 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V9_40Sx120_40V_120H

VIA V9_40Sx120_60V_120H
  LAYER m9 ;
    RECT -0.03 -0.084 0.03 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V9_40Sx120_60V_120H

VIA V9_40Sx120_80V_120H
  LAYER m9 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.06 0.058 0.06 ;
END V9_40Sx120_80V_120H

VIA V9_40Sx40_120H_40H
  LAYER m9 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v9 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m10 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V9_40Sx40_120H_40H

VIA V9_40Sx40_120V_40H
  LAYER m9 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v9 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m10 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V9_40Sx40_120V_40H

VIA V9_40Sx40_160H_40H
  LAYER m9 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v9 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m10 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V9_40Sx40_160H_40H

VIA V9_40Sx40_160V_40H
  LAYER m9 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v9 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m10 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V9_40Sx40_160V_40H

VIA V9_40Sx40_200H_40H
  LAYER m9 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v9 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m10 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V9_40Sx40_200H_40H

VIA V9_40Sx40_200V_40H
  LAYER m9 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v9 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m10 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V9_40Sx40_200V_40H

VIA V9_40Sx40_40V_40H
  LAYER m9 ;
    RECT -0.02 -0.044 0.02 0.044 ;
  LAYER v9 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m10 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V9_40Sx40_40V_40H

VIA V9_40Sx40_60V_40H
  LAYER m9 ;
    RECT -0.03 -0.044 0.03 0.044 ;
  LAYER v9 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m10 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V9_40Sx40_60V_40H

VIA V9_40Sx40_80H_40H
  LAYER m9 ;
    RECT -0.044 -0.04 0.044 0.04 ;
  LAYER v9 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m10 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V9_40Sx40_80H_40H

VIA V9_40Sx40_80V_40H
  LAYER m9 ;
    RECT -0.04 -0.044 0.04 0.044 ;
  LAYER v9 ;
    RECT -0.02 -0.02 0.02 0.02 ;
  LAYER m10 ;
    RECT -0.058 -0.02 0.058 0.02 ;
END V9_40Sx40_80V_40H

VIA V9_40Sx60_120H_60H
  LAYER m9 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v9 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m10 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V9_40Sx60_120H_60H

VIA V9_40Sx60_120V_60H
  LAYER m9 ;
    RECT -0.06 -0.054 0.06 0.054 ;
  LAYER v9 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m10 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V9_40Sx60_120V_60H

VIA V9_40Sx60_160H_60H
  LAYER m9 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v9 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m10 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V9_40Sx60_160H_60H

VIA V9_40Sx60_160V_60H
  LAYER m9 ;
    RECT -0.08 -0.054 0.08 0.054 ;
  LAYER v9 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m10 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V9_40Sx60_160V_60H

VIA V9_40Sx60_200H_60H
  LAYER m9 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v9 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m10 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V9_40Sx60_200H_60H

VIA V9_40Sx60_200V_60H
  LAYER m9 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v9 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m10 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V9_40Sx60_200V_60H

VIA V9_40Sx60_40V_60H
  LAYER m9 ;
    RECT -0.02 -0.054 0.02 0.054 ;
  LAYER v9 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m10 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V9_40Sx60_40V_60H

VIA V9_40Sx60_60V_60H
  LAYER m9 ;
    RECT -0.03 -0.054 0.03 0.054 ;
  LAYER v9 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m10 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V9_40Sx60_60V_60H

VIA V9_40Sx60_80H_60H
  LAYER m9 ;
    RECT -0.044 -0.04 0.044 0.04 ;
  LAYER v9 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m10 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V9_40Sx60_80H_60H

VIA V9_40Sx60_80V_60H
  LAYER m9 ;
    RECT -0.04 -0.054 0.04 0.054 ;
  LAYER v9 ;
    RECT -0.02 -0.03 0.02 0.03 ;
  LAYER m10 ;
    RECT -0.058 -0.03 0.058 0.03 ;
END V9_40Sx60_80V_60H

VIA V9_40Sx80_120H_80H
  LAYER m9 ;
    RECT -0.044 -0.06 0.044 0.06 ;
  LAYER v9 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m10 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V9_40Sx80_120H_80H

VIA V9_40Sx80_120V_80H
  LAYER m9 ;
    RECT -0.06 -0.064 0.06 0.064 ;
  LAYER v9 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m10 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V9_40Sx80_120V_80H

VIA V9_40Sx80_160H_80H
  LAYER m9 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v9 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m10 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V9_40Sx80_160H_80H

VIA V9_40Sx80_160V_80H
  LAYER m9 ;
    RECT -0.08 -0.064 0.08 0.064 ;
  LAYER v9 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m10 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V9_40Sx80_160V_80H

VIA V9_40Sx80_200H_80H
  LAYER m9 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v9 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m10 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V9_40Sx80_200H_80H

VIA V9_40Sx80_200V_80H
  LAYER m9 ;
    RECT -0.1 -0.064 0.1 0.064 ;
  LAYER v9 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m10 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V9_40Sx80_200V_80H

VIA V9_40Sx80_40V_80H
  LAYER m9 ;
    RECT -0.02 -0.064 0.02 0.064 ;
  LAYER v9 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m10 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V9_40Sx80_40V_80H

VIA V9_40Sx80_60V_80H
  LAYER m9 ;
    RECT -0.03 -0.064 0.03 0.064 ;
  LAYER v9 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m10 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V9_40Sx80_60V_80H

VIA V9_40Sx80_80H_80H
  LAYER m9 ;
    RECT -0.044 -0.04 0.044 0.04 ;
  LAYER v9 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m10 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V9_40Sx80_80H_80H

VIA V9_40Sx80_80V_80H
  LAYER m9 ;
    RECT -0.04 -0.064 0.04 0.064 ;
  LAYER v9 ;
    RECT -0.02 -0.04 0.02 0.04 ;
  LAYER m10 ;
    RECT -0.058 -0.04 0.058 0.04 ;
END V9_40Sx80_80V_80H

VIA V9_40x120_120V_120V
  LAYER m9 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V9_40x120_120V_120V

VIA V9_40x120_120V_160H
  LAYER m9 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V9_40x120_120V_160H

VIA V9_40x120_120V_160V
  LAYER m9 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V9_40x120_120V_160V

VIA V9_40x120_120V_200H
  LAYER m9 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V9_40x120_120V_200H

VIA V9_40x120_120V_200V
  LAYER m9 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V9_40x120_120V_200V

VIA V9_40x120_120V_80V
  LAYER m9 ;
    RECT -0.06 -0.084 0.06 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V9_40x120_120V_80V

VIA V9_40x120_160H_120V
  LAYER m9 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V9_40x120_160H_120V

VIA V9_40x120_160H_160H
  LAYER m9 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V9_40x120_160H_160H

VIA V9_40x120_160H_160V
  LAYER m9 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V9_40x120_160H_160V

VIA V9_40x120_160H_200H
  LAYER m9 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V9_40x120_160H_200H

VIA V9_40x120_160H_200V
  LAYER m9 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V9_40x120_160H_200V

VIA V9_40x120_160H_80V
  LAYER m9 ;
    RECT -0.044 -0.08 0.044 0.08 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V9_40x120_160H_80V

VIA V9_40x120_160V_120V
  LAYER m9 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V9_40x120_160V_120V

VIA V9_40x120_160V_160H
  LAYER m9 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V9_40x120_160V_160H

VIA V9_40x120_160V_160V
  LAYER m9 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V9_40x120_160V_160V

VIA V9_40x120_160V_200H
  LAYER m9 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V9_40x120_160V_200H

VIA V9_40x120_160V_200V
  LAYER m9 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V9_40x120_160V_200V

VIA V9_40x120_160V_80V
  LAYER m9 ;
    RECT -0.08 -0.084 0.08 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V9_40x120_160V_80V

VIA V9_40x120_200H_120V
  LAYER m9 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V9_40x120_200H_120V

VIA V9_40x120_200H_160H
  LAYER m9 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V9_40x120_200H_160H

VIA V9_40x120_200H_160V
  LAYER m9 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V9_40x120_200H_160V

VIA V9_40x120_200H_200H
  LAYER m9 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V9_40x120_200H_200H

VIA V9_40x120_200H_200V
  LAYER m9 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V9_40x120_200H_200V

VIA V9_40x120_200H_80V
  LAYER m9 ;
    RECT -0.044 -0.1 0.044 0.1 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V9_40x120_200H_80V

VIA V9_40x120_200V_120V
  LAYER m9 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V9_40x120_200V_120V

VIA V9_40x120_200V_160H
  LAYER m9 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V9_40x120_200V_160H

VIA V9_40x120_200V_160V
  LAYER m9 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V9_40x120_200V_160V

VIA V9_40x120_200V_200H
  LAYER m9 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V9_40x120_200V_200H

VIA V9_40x120_200V_200V
  LAYER m9 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V9_40x120_200V_200V

VIA V9_40x120_200V_80V
  LAYER m9 ;
    RECT -0.1 -0.084 0.1 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V9_40x120_200V_80V

VIA V9_40x120_80V_120V
  LAYER m9 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.06 -0.098 0.06 0.098 ;
END V9_40x120_80V_120V

VIA V9_40x120_80V_160H
  LAYER m9 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.08 0.058 0.08 ;
END V9_40x120_80V_160H

VIA V9_40x120_80V_160V
  LAYER m9 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.08 -0.098 0.08 0.098 ;
END V9_40x120_80V_160V

VIA V9_40x120_80V_200H
  LAYER m9 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.058 -0.1 0.058 0.1 ;
END V9_40x120_80V_200H

VIA V9_40x120_80V_200V
  LAYER m9 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.1 -0.098 0.1 0.098 ;
END V9_40x120_80V_200V

VIA V9_40x120_80V_80V
  LAYER m9 ;
    RECT -0.04 -0.084 0.04 0.084 ;
  LAYER v9 ;
    RECT -0.02 -0.06 0.02 0.06 ;
  LAYER m10 ;
    RECT -0.04 -0.098 0.04 0.098 ;
END V9_40x120_80V_80V

VIA V9_60Sx40_120H_40H
  LAYER m9 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v9 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m10 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V9_60Sx40_120H_40H

VIA V9_60Sx40_120V_40H
  LAYER m9 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v9 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m10 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V9_60Sx40_120V_40H

VIA V9_60Sx40_160H_40H
  LAYER m9 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v9 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m10 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V9_60Sx40_160H_40H

VIA V9_60Sx40_160V_40H
  LAYER m9 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v9 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m10 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V9_60Sx40_160V_40H

VIA V9_60Sx40_200H_40H
  LAYER m9 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v9 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m10 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V9_60Sx40_200H_40H

VIA V9_60Sx40_200V_40H
  LAYER m9 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v9 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m10 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V9_60Sx40_200V_40H

VIA V9_60Sx40_60V_40H
  LAYER m9 ;
    RECT -0.03 -0.044 0.03 0.044 ;
  LAYER v9 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m10 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V9_60Sx40_60V_40H

VIA V9_60Sx40_80H_40H
  LAYER m9 ;
    RECT -0.054 -0.04 0.054 0.04 ;
  LAYER v9 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m10 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V9_60Sx40_80H_40H

VIA V9_60Sx40_80V_40H
  LAYER m9 ;
    RECT -0.04 -0.044 0.04 0.044 ;
  LAYER v9 ;
    RECT -0.03 -0.02 0.03 0.02 ;
  LAYER m10 ;
    RECT -0.068 -0.02 0.068 0.02 ;
END V9_60Sx40_80V_40H

VIA V9_60Sx60_120H_60H
  LAYER m9 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v9 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m10 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V9_60Sx60_120H_60H

VIA V9_60Sx60_120V_60H
  LAYER m9 ;
    RECT -0.06 -0.054 0.06 0.054 ;
  LAYER v9 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m10 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V9_60Sx60_120V_60H

VIA V9_60Sx60_160H_60H
  LAYER m9 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v9 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m10 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V9_60Sx60_160H_60H

VIA V9_60Sx60_160V_60H
  LAYER m9 ;
    RECT -0.08 -0.054 0.08 0.054 ;
  LAYER v9 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m10 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V9_60Sx60_160V_60H

VIA V9_60Sx60_200H_60H
  LAYER m9 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v9 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m10 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V9_60Sx60_200H_60H

VIA V9_60Sx60_200V_60H
  LAYER m9 ;
    RECT -0.1 -0.054 0.1 0.054 ;
  LAYER v9 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m10 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V9_60Sx60_200V_60H

VIA V9_60Sx60_60V_60H
  LAYER m9 ;
    RECT -0.03 -0.054 0.03 0.054 ;
  LAYER v9 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m10 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V9_60Sx60_60V_60H

VIA V9_60Sx60_80H_60H
  LAYER m9 ;
    RECT -0.054 -0.04 0.054 0.04 ;
  LAYER v9 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m10 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V9_60Sx60_80H_60H

VIA V9_60Sx60_80V_60H
  LAYER m9 ;
    RECT -0.04 -0.054 0.04 0.054 ;
  LAYER v9 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER m10 ;
    RECT -0.068 -0.03 0.068 0.03 ;
END V9_60Sx60_80V_60H

VIA V9_60Sx80_120H_80H
  LAYER m9 ;
    RECT -0.054 -0.06 0.054 0.06 ;
  LAYER v9 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m10 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V9_60Sx80_120H_80H

VIA V9_60Sx80_120V_80H
  LAYER m9 ;
    RECT -0.06 -0.064 0.06 0.064 ;
  LAYER v9 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m10 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V9_60Sx80_120V_80H

VIA V9_60Sx80_160H_80H
  LAYER m9 ;
    RECT -0.054 -0.08 0.054 0.08 ;
  LAYER v9 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m10 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V9_60Sx80_160H_80H

VIA V9_60Sx80_160V_80H
  LAYER m9 ;
    RECT -0.08 -0.064 0.08 0.064 ;
  LAYER v9 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m10 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V9_60Sx80_160V_80H

VIA V9_60Sx80_200H_80H
  LAYER m9 ;
    RECT -0.054 -0.1 0.054 0.1 ;
  LAYER v9 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m10 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V9_60Sx80_200H_80H

VIA V9_60Sx80_200V_80H
  LAYER m9 ;
    RECT -0.1 -0.064 0.1 0.064 ;
  LAYER v9 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m10 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V9_60Sx80_200V_80H

VIA V9_60Sx80_60V_80H
  LAYER m9 ;
    RECT -0.03 -0.064 0.03 0.064 ;
  LAYER v9 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m10 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V9_60Sx80_60V_80H

VIA V9_60Sx80_80H_80H
  LAYER m9 ;
    RECT -0.054 -0.04 0.054 0.04 ;
  LAYER v9 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m10 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V9_60Sx80_80H_80H

VIA V9_60Sx80_80V_80H
  LAYER m9 ;
    RECT -0.04 -0.064 0.04 0.064 ;
  LAYER v9 ;
    RECT -0.03 -0.04 0.03 0.04 ;
  LAYER m10 ;
    RECT -0.068 -0.04 0.068 0.04 ;
END V9_60Sx80_80V_80H

VIA V9_80x40S_120H_80V
  LAYER m9 ;
    RECT -0.064 -0.06 0.064 0.06 ;
  LAYER v9 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m10 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V9_80x40S_120H_80V

VIA V9_80x40S_120V_80V
  LAYER m9 ;
    RECT -0.06 -0.044 0.06 0.044 ;
  LAYER v9 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m10 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V9_80x40S_120V_80V

VIA V9_80x40S_160H_80V
  LAYER m9 ;
    RECT -0.064 -0.08 0.064 0.08 ;
  LAYER v9 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m10 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V9_80x40S_160H_80V

VIA V9_80x40S_160V_80V
  LAYER m9 ;
    RECT -0.08 -0.044 0.08 0.044 ;
  LAYER v9 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m10 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V9_80x40S_160V_80V

VIA V9_80x40S_200H_80V
  LAYER m9 ;
    RECT -0.064 -0.1 0.064 0.1 ;
  LAYER v9 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m10 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V9_80x40S_200H_80V

VIA V9_80x40S_200V_80V
  LAYER m9 ;
    RECT -0.1 -0.044 0.1 0.044 ;
  LAYER v9 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m10 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V9_80x40S_200V_80V

VIA V9_80x40S_80H_80V
  LAYER m9 ;
    RECT -0.064 -0.04 0.064 0.04 ;
  LAYER v9 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m10 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V9_80x40S_80H_80V

VIA V9_80x40S_80V_80V
  LAYER m9 ;
    RECT -0.04 -0.044 0.04 0.044 ;
  LAYER v9 ;
    RECT -0.04 -0.02 0.04 0.02 ;
  LAYER m10 ;
    RECT -0.04 -0.058 0.04 0.058 ;
END V9_80x40S_80V_80V

VIA VG_DUMMY
  LAYER bm0 ;
    RECT -0.01 -0.007 0.01 0.007 ;
  LAYER vg ;
    RECT -0.01 -0.007 0.01 0.007 ;
  LAYER m0 ;
    RECT -0.01 -0.007 0.01 0.007 ;
END VG_DUMMY

NONDEFAULTRULE ndr_defaultW_3T_noSh
  HARDSPACING ;
  LAYER bsb
    WIDTH 32 ;
    SPACING 0.001 ;
  END bsb
  LAYER bm5
    WIDTH 2 ;
    SPACING 2 ;
  END bm5
  LAYER bm4
    WIDTH 0.54 ;
    SPACING 0.54 ;
  END bm4
  LAYER bm3
    WIDTH 0.54 ;
    SPACING 0.54 ;
  END bm3
  LAYER bm2
    WIDTH 0.24 ;
    SPACING 0.14 ;
  END bm2
  LAYER bm1
    WIDTH 0.16 ;
    SPACING 0.14 ;
  END bm1
  LAYER bm0
    WIDTH 0.08 ;
    SPACING 0.08 ;
  END bm0
  LAYER m0
    WIDTH 0.02 ;
    SPACING 0.016 ;
  END m0
  LAYER m1
    WIDTH 0.03 ;
    SPACING 0.02 ;
  END m1
  LAYER m2
    WIDTH 0.02 ;
    SPACING 0.016 ;
  END m2
  LAYER m3
    WIDTH 0.024 ;
    SPACING 0.016 ;
  END m3
  LAYER m4
    WIDTH 0.024 ;
    SPACING 0.016 ;
  END m4
  LAYER m5
    WIDTH 0.04 ;
    SPACING 0.08 ;
  END m5
  LAYER m6
    WIDTH 0.04 ;
    SPACING 0.08 ;
  END m6
  LAYER m7
    WIDTH 0.04 ;
    SPACING 0.08 ;
  END m7
  LAYER m8
    WIDTH 0.04 ;
    SPACING 0.08 ;
  END m8
  LAYER m9
    WIDTH 0.04 ;
    SPACING 0.08 ;
  END m9
  LAYER m10
    WIDTH 0.04 ;
    SPACING 0.08 ;
  END m10
  LAYER m11
    WIDTH 0.06 ;
    SPACING 0.12 ;
  END m11
  LAYER m12
    WIDTH 0.06 ;
    SPACING 0.12 ;
  END m12
  LAYER m13
    WIDTH 0.08 ;
    SPACING 0.16 ;
  END m13
  LAYER m14
    WIDTH 0.08 ;
    SPACING 0.16 ;
  END m14
END ndr_defaultW_3T_noSh

NONDEFAULTRULE ndr_defaultW_3T_Sh
  HARDSPACING ;
  LAYER bsb
    WIDTH 32 ;
    SPACING 0.001 ;
  END bsb
  LAYER bm5
    WIDTH 2 ;
    SPACING 2 ;
  END bm5
  LAYER bm4
    WIDTH 0.54 ;
    SPACING 0.54 ;
  END bm4
  LAYER bm3
    WIDTH 0.54 ;
    SPACING 0.54 ;
  END bm3
  LAYER bm2
    WIDTH 0.24 ;
    SPACING 0.14 ;
  END bm2
  LAYER bm1
    WIDTH 0.16 ;
    SPACING 0.14 ;
  END bm1
  LAYER bm0
    WIDTH 0.08 ;
    SPACING 0.08 ;
  END bm0
  LAYER m0
    WIDTH 0.02 ;
    SPACING 0.016 ;
  END m0
  LAYER m1
    WIDTH 0.03 ;
    SPACING 0.02 ;
  END m1
  LAYER m2
    WIDTH 0.02 ;
    SPACING 0.016 ;
  END m2
  LAYER m3
    WIDTH 0.024 ;
    SPACING 0.016 ;
  END m3
  LAYER m4
    WIDTH 0.024 ;
    SPACING 0.016 ;
  END m4
  LAYER m5
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m5
  LAYER m6
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m6
  LAYER m7
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m7
  LAYER m8
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m8
  LAYER m9
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m9
  LAYER m10
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m10
  LAYER m11
    WIDTH 0.06 ;
    SPACING 0.06 ;
  END m11
  LAYER m12
    WIDTH 0.06 ;
    SPACING 0.06 ;
  END m12
  LAYER m13
    WIDTH 0.08 ;
    SPACING 0.08 ;
  END m13
  LAYER m14
    WIDTH 0.08 ;
    SPACING 0.08 ;
  END m14
END ndr_defaultW_3T_Sh

NONDEFAULTRULE ndr_wide_wire_pat_80
  HARDSPACING ;
  LAYER bsb
    WIDTH 32 ;
    SPACING 0.001 ;
  END bsb
  LAYER bm5
    WIDTH 2 ;
    SPACING 2 ;
  END bm5
  LAYER bm4
    WIDTH 0.54 ;
    SPACING 0.54 ;
  END bm4
  LAYER bm3
    WIDTH 0.54 ;
    SPACING 0.54 ;
  END bm3
  LAYER bm2
    WIDTH 0.24 ;
    SPACING 0.14 ;
  END bm2
  LAYER bm1
    WIDTH 0.16 ;
    SPACING 0.14 ;
  END bm1
  LAYER bm0
    WIDTH 0.08 ;
    SPACING 0.08 ;
  END bm0
  LAYER m0
    WIDTH 0.02 ;
    SPACING 0.016 ;
  END m0
  LAYER m1
    WIDTH 0.03 ;
    SPACING 0.02 ;
  END m1
  LAYER m2
    WIDTH 0.02 ;
    SPACING 0.016 ;
  END m2
  LAYER m3
    WIDTH 0.044 ;
    SPACING 0.016 ;
  END m3
  LAYER m4
    WIDTH 0.044 ;
    SPACING 0.016 ;
  END m4
  LAYER m5
    WIDTH 0.08 ;
    SPACING 0.04 ;
  END m5
  LAYER m6
    WIDTH 0.08 ;
    SPACING 0.04 ;
  END m6
  LAYER m7
    WIDTH 0.08 ;
    SPACING 0.04 ;
  END m7
  LAYER m8
    WIDTH 0.08 ;
    SPACING 0.04 ;
  END m8
  LAYER m9
    WIDTH 0.08 ;
    SPACING 0.04 ;
  END m9
  LAYER m10
    WIDTH 0.08 ;
    SPACING 0.04 ;
  END m10
  LAYER m11
    WIDTH 0.12 ;
    SPACING 0.06 ;
  END m11
  LAYER m12
    WIDTH 0.12 ;
    SPACING 0.06 ;
  END m12
  LAYER m13
    WIDTH 0.16 ;
    SPACING 0.08 ;
  END m13
  LAYER m14
    WIDTH 0.16 ;
    SPACING 0.08 ;
  END m14
END ndr_wide_wire_pat_80

NONDEFAULTRULE ndr_wide_wire_pat_160
  HARDSPACING ;
  LAYER bsb
    WIDTH 32 ;
    SPACING 0.001 ;
  END bsb
  LAYER bm5
    WIDTH 2 ;
    SPACING 2 ;
  END bm5
  LAYER bm4
    WIDTH 0.54 ;
    SPACING 0.54 ;
  END bm4
  LAYER bm3
    WIDTH 0.54 ;
    SPACING 0.54 ;
  END bm3
  LAYER bm2
    WIDTH 0.24 ;
    SPACING 0.14 ;
  END bm2
  LAYER bm1
    WIDTH 0.16 ;
    SPACING 0.14 ;
  END bm1
  LAYER bm0
    WIDTH 0.08 ;
    SPACING 0.08 ;
  END bm0
  LAYER m0
    WIDTH 0.02 ;
    SPACING 0.016 ;
  END m0
  LAYER m1
    WIDTH 0.03 ;
    SPACING 0.02 ;
  END m1
  LAYER m2
    WIDTH 0.02 ;
    SPACING 0.016 ;
  END m2
  LAYER m3
    WIDTH 0.044 ;
    SPACING 0.016 ;
  END m3
  LAYER m4
    WIDTH 0.044 ;
    SPACING 0.016 ;
  END m4
  LAYER m5
    WIDTH 0.16 ;
    SPACING 0.04 ;
  END m5
  LAYER m6
    WIDTH 0.16 ;
    SPACING 0.04 ;
  END m6
  LAYER m7
    WIDTH 0.16 ;
    SPACING 0.04 ;
  END m7
  LAYER m8
    WIDTH 0.16 ;
    SPACING 0.04 ;
  END m8
  LAYER m9
    WIDTH 0.16 ;
    SPACING 0.04 ;
  END m9
  LAYER m10
    WIDTH 0.16 ;
    SPACING 0.04 ;
  END m10
  LAYER m11
    WIDTH 0.24 ;
    SPACING 0.06 ;
  END m11
  LAYER m12
    WIDTH 0.24 ;
    SPACING 0.06 ;
  END m12
  LAYER m13
    WIDTH 0.32 ;
    SPACING 0.08 ;
  END m13
  LAYER m14
    WIDTH 0.32 ;
    SPACING 0.08 ;
  END m14
END ndr_wide_wire_pat_160

NONDEFAULTRULE ndr_2W_StrongSh
  HARDSPACING ;
  LAYER bsb
    WIDTH 32 ;
    SPACING 0.001 ;
  END bsb
  LAYER bm5
    WIDTH 2 ;
    SPACING 2 ;
  END bm5
  LAYER bm4
    WIDTH 0.54 ;
    SPACING 0.54 ;
  END bm4
  LAYER bm3
    WIDTH 0.54 ;
    SPACING 0.54 ;
  END bm3
  LAYER bm2
    WIDTH 0.24 ;
    SPACING 0.14 ;
  END bm2
  LAYER bm1
    WIDTH 0.16 ;
    SPACING 0.14 ;
  END bm1
  LAYER bm0
    WIDTH 0.08 ;
    SPACING 0.08 ;
  END bm0
  LAYER m0
    WIDTH 0.02 ;
    SPACING 0.016 ;
  END m0
  LAYER m1
    WIDTH 0.03 ;
    SPACING 0.02 ;
  END m1
  LAYER m2
    WIDTH 0.02 ;
    SPACING 0.016 ;
  END m2
  LAYER m3
    WIDTH 0.024 ;
    SPACING 0.016 ;
  END m3
  LAYER m4
    WIDTH 0.024 ;
    SPACING 0.016 ;
  END m4
  LAYER m5
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m5
  LAYER m6
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m6
  LAYER m7
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m7
  LAYER m8
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m8
  LAYER m9
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m9
  LAYER m10
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m10
  LAYER m11
    WIDTH 0.06 ;
    SPACING 0.06 ;
  END m11
  LAYER m12
    WIDTH 0.06 ;
    SPACING 0.06 ;
  END m12
  LAYER m13
    WIDTH 0.16 ;
    SPACING 0.08 ;
  END m13
  LAYER m14
    WIDTH 0.16 ;
    SPACING 0.08 ;
  END m14
END ndr_2W_StrongSh

NONDEFAULTRULE rm_leaf
  HARDSPACING ;
  LAYER bsb
    WIDTH 32 ;
    SPACING 0.001 ;
  END bsb
  LAYER bm5
    WIDTH 2 ;
    SPACING 2 ;
  END bm5
  LAYER bm4
    WIDTH 0.54 ;
    SPACING 0.54 ;
  END bm4
  LAYER bm3
    WIDTH 0.54 ;
    SPACING 0.54 ;
  END bm3
  LAYER bm2
    WIDTH 0.24 ;
    SPACING 0.14 ;
  END bm2
  LAYER bm1
    WIDTH 0.16 ;
    SPACING 0.14 ;
  END bm1
  LAYER bm0
    WIDTH 0.08 ;
    SPACING 0.08 ;
  END bm0
  LAYER m0
    WIDTH 0.02 ;
    SPACING 0.016 ;
  END m0
  LAYER m1
    WIDTH 0.03 ;
    SPACING 0.02 ;
  END m1
  LAYER m2
    WIDTH 0.02 ;
    SPACING 0.016 ;
  END m2
  LAYER m3
    WIDTH 0.024 ;
    SPACING 0.016 ;
  END m3
  LAYER m4
    WIDTH 0.024 ;
    SPACING 0.016 ;
  END m4
  LAYER m5
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m5
  LAYER m6
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m6
  LAYER m7
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m7
  LAYER m8
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m8
  LAYER m9
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m9
  LAYER m10
    WIDTH 0.04 ;
    SPACING 0.04 ;
  END m10
  LAYER m11
    WIDTH 0.06 ;
    SPACING 0.06 ;
  END m11
  LAYER m12
    WIDTH 0.06 ;
    SPACING 0.06 ;
  END m12
  LAYER m13
    WIDTH 0.08 ;
    SPACING 0.08 ;
  END m13
  LAYER m14
    WIDTH 0.08 ;
    SPACING 0.08 ;
  END m14
END rm_leaf

SITE unit_100
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.1 BY 0.27 ;
END unit_100

SITE core_100
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.1 BY 0.27 ;
END core_100

SITE core2h_100
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.1 BY 0.54 ;
END core2h_100

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.05 BY 0.18 ;
END unit

SITE core
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.05 BY 0.18 ;
END core

SITE bonuscore
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.25 BY 0.18 ;
END bonuscore

SITE core2h
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.05 BY 0.36 ;
END core2h

SITE core4h
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.05 BY 0.72 ;
END core4h

MACRO i0maoi222aa1n02x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.4 BY 0.18 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m0 ;
        RECT 0.283 0.062 0.392 0.082 ;
      LAYER vg ;
        RECT 0.293 0.062 0.307 0.082 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.001288 ;
  END a
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m0 ;
        RECT 0.308 0.026 0.392 0.046 ;
      LAYER vg ;
        RECT 0.343 0.026 0.357 0.046 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.001288 ;
  END b
  PIN c
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m0 ;
        RECT 0.058 0.062 0.167 0.082 ;
      LAYER vg ;
        RECT 0.143 0.062 0.157 0.082 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.001288 ;
  END c
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m1 ;
        RECT 0.21 0.015 0.24 0.093 ;
      LAYER m0 ;
        RECT 0.183 0.062 0.242 0.082 ;
      LAYER v0 ;
        RECT 0.21 0.062 0.24 0.082 ;
      LAYER vg ;
        RECT 0.193 0.062 0.207 0.082 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.001288 ;
  END d
  PIN e
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m0 ;
        RECT 0.058 0.134 0.142 0.154 ;
      LAYER vg ;
        RECT 0.093 0.134 0.107 0.154 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.001288 ;
  END e
  PIN f
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m0 ;
        RECT 0.008 0.026 0.092 0.046 ;
      LAYER vg ;
        RECT 0.043 0.026 0.057 0.046 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.001288 ;
  END f
  PIN o1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m1 ;
        RECT 0.26 0.015 0.29 0.129 ;
      LAYER m0 ;
        RECT 0.108 0.026 0.292 0.046 ;
        RECT 0.258 0.098 0.342 0.118 ;
      LAYER v0 ;
        RECT 0.26 0.026 0.29 0.046 ;
        RECT 0.26 0.098 0.29 0.118 ;
      LAYER vt ;
        RECT 0.117 0.026 0.133 0.046 ;
        RECT 0.267 0.026 0.283 0.046 ;
        RECT 0.317 0.098 0.333 0.118 ;
    END
    ANTENNADIFFAREA 0.004968 ;
  END o1
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER bm0 ;
        RECT -0.085 0.14 0.485 0.22 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER bm0 ;
        RECT -0.085 -0.04 0.485 0.04 ;
    END
  END vssx
  OBS
    LAYER m0 ;
      RECT 0.158 0.134 0.392 0.154 ;
      RECT 0.258 0.098 0.342 0.118 ;
      RECT 0.008 0.098 0.242 0.118 ;
      RECT 0.183 0.062 0.242 0.082 ;
      RECT 0.108 0.026 0.292 0.046 ;
      RECT 0.158 0.134 0.392 0.154 ;
      RECT 0.008 0.098 0.242 0.118 ;
    LAYER dvb ;
      RECT -0.0655 0.171 0.4655 0.189 ;
      RECT -0.0655 -0.009 0.4655 0.009 ;
    LAYER ndiff ;
      RECT 0.257 0.028 0.393 0.074 ;
      RECT 0.007 0.028 0.243 0.074 ;
    LAYER pdiff ;
      RECT 0.257 0.106 0.393 0.152 ;
      RECT 0.007 0.106 0.243 0.152 ;
    LAYER tcn ;
      RECT 0.067 0.098 0.083 0.187 ;
      RECT 0.367 0.098 0.383 0.157 ;
      RECT 0.317 0.098 0.333 0.157 ;
      RECT 0.267 0.098 0.283 0.157 ;
      RECT 0.217 0.098 0.233 0.157 ;
      RECT 0.167 0.098 0.183 0.157 ;
      RECT 0.117 0.098 0.133 0.157 ;
      RECT 0.017 0.098 0.033 0.157 ;
      RECT 0.367 -0.007 0.383 0.082 ;
      RECT 0.317 0.023 0.333 0.082 ;
      RECT 0.267 0.023 0.283 0.082 ;
      RECT 0.217 -0.007 0.233 0.082 ;
      RECT 0.167 0.023 0.183 0.082 ;
      RECT 0.117 0.023 0.133 0.082 ;
      RECT 0.067 0.023 0.083 0.082 ;
      RECT 0.017 -0.007 0.033 0.082 ;
    LAYER devflav_n5_id ;
      RECT 0 0 0.4 0.09 ;
    LAYER devflav_p5_id ;
      RECT 0 0.09 0.4 0.18 ;
  END
END i0maoi222aa1n02x5

MACRO i0mbff000aa1n30x5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.85 BY 0.18 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m0 ;
        RECT 0.033 0.026 0.317 0.046 ;
      LAYER vg ;
        RECT 0.043 0.026 0.057 0.046 ;
        RECT 0.093 0.026 0.107 0.046 ;
        RECT 0.193 0.026 0.207 0.046 ;
        RECT 0.243 0.026 0.257 0.046 ;
        RECT 0.293 0.026 0.307 0.046 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.00784 ;
  END a
  PIN o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m1 ;
        RECT 0.36 0.015 0.39 0.093 ;
        RECT 0.46 0.015 0.49 0.093 ;
        RECT 0.56 0.015 0.59 0.093 ;
        RECT 0.66 0.015 0.69 0.093 ;
        RECT 0.76 0.015 0.79 0.093 ;
      LAYER m0 ;
        RECT 0.358 0.026 0.792 0.082 ;
      LAYER vt ;
        RECT 0.367 0.026 0.383 0.082 ;
        RECT 0.467 0.026 0.483 0.082 ;
        RECT 0.567 0.026 0.583 0.082 ;
        RECT 0.667 0.026 0.683 0.082 ;
        RECT 0.767 0.026 0.783 0.082 ;
      LAYER v0 ;
        RECT 0.36 0.026 0.39 0.082 ;
        RECT 0.46 0.026 0.49 0.082 ;
        RECT 0.56 0.026 0.59 0.082 ;
        RECT 0.66 0.026 0.69 0.082 ;
        RECT 0.76 0.026 0.79 0.082 ;
    END
    PROPERTY LEF58_MUSTJOINALLPORTS "MUSTJOINALLPORTS ;" ;
    ANTENNADIFFAREA 0.02016 ;
  END o
  PIN vcc
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER bm0 ;
        RECT -0.085 0.14 0.935 0.22 ;
    END
  END vcc
  PIN vssx
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER bm0 ;
        RECT -0.085 -0.04 0.935 0.04 ;
    END
  END vssx
  OBS
    LAYER m0 ;
      RECT 0.058 0.134 0.817 0.154 ;
      RECT 0.358 0.026 0.792 0.082 ;
    LAYER vg ;
      RECT 0.793 0.134 0.807 0.154 ;
      RECT 0.743 0.134 0.757 0.154 ;
      RECT 0.693 0.134 0.707 0.154 ;
      RECT 0.643 0.134 0.657 0.154 ;
      RECT 0.593 0.134 0.607 0.154 ;
      RECT 0.543 0.134 0.557 0.154 ;
      RECT 0.493 0.134 0.507 0.154 ;
      RECT 0.443 0.134 0.457 0.154 ;
      RECT 0.393 0.134 0.407 0.154 ;
      RECT 0.343 0.134 0.357 0.154 ;
    LAYER m0 ;
      RECT 0.058 0.134 0.817 0.154 ;
    LAYER dvb ;
      RECT -0.0655 0.171 0.9155 0.189 ;
      RECT -0.0655 -0.009 0.9155 0.009 ;
    LAYER ndiff ;
      RECT 0.157 0.023 0.843 0.079 ;
      RECT 0.007 0.023 0.143 0.079 ;
    LAYER pdiff ;
      RECT 0.157 0.101 0.843 0.157 ;
      RECT 0.007 0.101 0.143 0.157 ;
    LAYER tcn ;
      RECT 0.817 0.098 0.833 0.187 ;
      RECT 0.717 0.098 0.733 0.187 ;
      RECT 0.617 0.098 0.633 0.187 ;
      RECT 0.517 0.098 0.533 0.187 ;
      RECT 0.417 0.098 0.433 0.187 ;
      RECT 0.317 0.098 0.333 0.187 ;
      RECT 0.217 0.098 0.233 0.187 ;
      RECT 0.117 0.098 0.133 0.187 ;
      RECT 0.017 0.098 0.033 0.187 ;
      RECT 0.767 0.023 0.783 0.157 ;
      RECT 0.667 0.023 0.683 0.157 ;
      RECT 0.567 0.023 0.583 0.157 ;
      RECT 0.467 0.023 0.483 0.157 ;
      RECT 0.367 0.023 0.383 0.157 ;
      RECT 0.267 0.023 0.283 0.157 ;
      RECT 0.167 0.023 0.183 0.157 ;
      RECT 0.067 0.023 0.083 0.157 ;
      RECT 0.817 -0.007 0.833 0.082 ;
      RECT 0.717 -0.007 0.733 0.082 ;
      RECT 0.617 -0.007 0.633 0.082 ;
      RECT 0.517 -0.007 0.533 0.082 ;
      RECT 0.417 -0.007 0.433 0.082 ;
      RECT 0.317 -0.007 0.333 0.082 ;
      RECT 0.217 -0.007 0.233 0.082 ;
      RECT 0.117 -0.007 0.133 0.082 ;
      RECT 0.017 -0.007 0.033 0.082 ;
    LAYER devflav_n5_id ;
      RECT 0 0 0.85 0.09 ;
    LAYER devflav_p5_id ;
      RECT 0 0.09 0.85 0.18 ;
  END
END i0mbff000aa1n30x5

MACRO i0mzh50basetbe04x
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  SIZE 0.05 BY 0.18 ;
  SYMMETRY X Y ;
  SITE core ;
END i0mzh50basetbe04x

MACRO i0mzh50baseysx04x
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  SIZE 0.2 BY 0.18 ;
  SYMMETRY X Y ;
  SITE core ;
END i0mzh50baseysx04x

MACRO i0mzh50basecxe04x
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  SIZE 0.2 BY 0.18 ;
  SYMMETRY X Y ;
  SITE core ;
END i0mzh50basecxe04x

END LIBRARY
